module half_adder(S, Cout, A, B);
    input A, B;
    output S, Cout;

    assign S = A ^ B;
    assign Cout = A & B;

endmodule