module not_(data_result, data_operandA);

    input [31:0] data_operandA;
    output [31:0] data_result;
    
    not NOT0(data_result[0], data_operandA[0]);
    not NOT1(data_result[1], data_operandA[1]);
    not NOT2(data_result[2], data_operandA[2]);
    not NOT3(data_result[3], data_operandA[3]);
    not NOT4(data_result[4], data_operandA[4]);
    not NOT5(data_result[5], data_operandA[5]);
    not NOT6(data_result[6], data_operandA[6]);
    not NOT7(data_result[7], data_operandA[7]);
    not NOT8(data_result[8], data_operandA[8]);
    not NOT9(data_result[9], data_operandA[9]);
    not NOT10(data_result[10], data_operandA[10]);
    not NOT11(data_result[11], data_operandA[11]);
    not NOT12(data_result[12], data_operandA[12]);
    not NOT13(data_result[13], data_operandA[13]);
    not NOT14(data_result[14], data_operandA[14]);
    not NOT15(data_result[15], data_operandA[15]);
    not NOT16(data_result[16], data_operandA[16]);
    not NOT17(data_result[17], data_operandA[17]);
    not NOT18(data_result[18], data_operandA[18]);
    not NOT19(data_result[19], data_operandA[19]);
    not NOT20(data_result[20], data_operandA[20]);
    not NOT21(data_result[21], data_operandA[21]);
    not NOT22(data_result[22], data_operandA[22]);
    not NOT23(data_result[23], data_operandA[23]);
    not NOT24(data_result[24], data_operandA[24]);
    not NOT25(data_result[25], data_operandA[25]);
    not NOT26(data_result[26], data_operandA[26]);
    not NOT27(data_result[27], data_operandA[27]);
    not NOT28(data_result[28], data_operandA[28]);
    not NOT29(data_result[29], data_operandA[29]);
    not NOT30(data_result[30], data_operandA[30]);
    not NOT31(data_result[31], data_operandA[31]);
endmodule