module wallacetree_32(Pout, Cout, A, B, C, ctrl_MULT, clock, ready);
    input [31:0] A, B;
    input C, ctrl_MULT, clock;
    output [31:0] Pout;
    output ready, Cout;

    wire [63:0] P;

    // all ANDs

    wire zero;
    assign zero = 1'b0;

    //level 1
    wire AND_A0_B0;
    and and_a0_b0(AND_A0_B0, A[0], B[0]);
    wire P_A0_B0, Cout_A0_B0;
    half_adder add_a0_b0(P_A0_B0, Cout_A0_B0, zero, AND_A0_B0);

    wire AND_A1_B0;
    and and_a1_b0(AND_A1_B0, A[1], B[0]);
    wire P_A1_B0, Cout_A1_B0;
    half_adder add_a1_b0(P_A1_B0, Cout_A1_B0, zero, AND_A1_B0);

    wire AND_A2_B0;
    and and_a2_b0(AND_A2_B0, A[2], B[0]);
    wire P_A2_B0, Cout_A2_B0;
    half_adder add_a2_b0(P_A2_B0, Cout_A2_B0, zero, AND_A2_B0);

    wire AND_A3_B0;
    and and_a3_b0(AND_A3_B0, A[3], B[0]);
    wire P_A3_B0, Cout_A3_B0;
    half_adder add_a3_b0(P_A3_B0, Cout_A3_B0, zero, AND_A3_B0);

    wire AND_A4_B0;
    and and_a4_b0(AND_A4_B0, A[4], B[0]);
    wire P_A4_B0, Cout_A4_B0;
    half_adder add_a4_b0(P_A4_B0, Cout_A4_B0, zero, AND_A4_B0);

    wire AND_A5_B0;
    and and_a5_b0(AND_A5_B0, A[5], B[0]);
    wire P_A5_B0, Cout_A5_B0;
    half_adder add_a5_b0(P_A5_B0, Cout_A5_B0, zero, AND_A5_B0);

    wire AND_A6_B0;
    and and_a6_b0(AND_A6_B0, A[6], B[0]);
    wire P_A6_B0, Cout_A6_B0;
    half_adder add_a6_b0(P_A6_B0, Cout_A6_B0, zero, AND_A6_B0);

    wire AND_A7_B0;
    and and_a7_b0(AND_A7_B0, A[7], B[0]);
    wire P_A7_B0, Cout_A7_B0;
    half_adder add_a7_b0(P_A7_B0, Cout_A7_B0, zero, AND_A7_B0);

    wire AND_A8_B0;
    and and_a8_b0(AND_A8_B0, A[8], B[0]);
    wire P_A8_B0, Cout_A8_B0;
    half_adder add_a8_b0(P_A8_B0, Cout_A8_B0, zero, AND_A8_B0);

    wire AND_A9_B0;
    and and_a9_b0(AND_A9_B0, A[9], B[0]);
    wire P_A9_B0, Cout_A9_B0;
    half_adder add_a9_b0(P_A9_B0, Cout_A9_B0, zero, AND_A9_B0);

    wire AND_A10_B0;
    and and_a10_b0(AND_A10_B0, A[10], B[0]);
    wire P_A10_B0, Cout_A10_B0;
    half_adder add_a10_b0(P_A10_B0, Cout_A10_B0, zero, AND_A10_B0);

    wire AND_A11_B0;
    and and_a11_b0(AND_A11_B0, A[11], B[0]);
    wire P_A11_B0, Cout_A11_B0;
    half_adder add_a11_b0(P_A11_B0, Cout_A11_B0, zero, AND_A11_B0);

    wire AND_A12_B0;
    and and_a12_b0(AND_A12_B0, A[12], B[0]);
    wire P_A12_B0, Cout_A12_B0;
    half_adder add_a12_b0(P_A12_B0, Cout_A12_B0, zero, AND_A12_B0);

    wire AND_A13_B0;
    and and_a13_b0(AND_A13_B0, A[13], B[0]);
    wire P_A13_B0, Cout_A13_B0;
    half_adder add_a13_b0(P_A13_B0, Cout_A13_B0, zero, AND_A13_B0);

    wire AND_A14_B0;
    and and_a14_b0(AND_A14_B0, A[14], B[0]);
    wire P_A14_B0, Cout_A14_B0;
    half_adder add_a14_b0(P_A14_B0, Cout_A14_B0, zero, AND_A14_B0);

    wire AND_A15_B0;
    and and_a15_b0(AND_A15_B0, A[15], B[0]);
    wire P_A15_B0, Cout_A15_B0;
    half_adder add_a15_b0(P_A15_B0, Cout_A15_B0, zero, AND_A15_B0);

    wire AND_A16_B0;
    and and_a16_b0(AND_A16_B0, A[16], B[0]);
    wire P_A16_B0, Cout_A16_B0;
    half_adder add_a16_b0(P_A16_B0, Cout_A16_B0, zero, AND_A16_B0);

    wire AND_A17_B0;
    and and_a17_b0(AND_A17_B0, A[17], B[0]);
    wire P_A17_B0, Cout_A17_B0;
    half_adder add_a17_b0(P_A17_B0, Cout_A17_B0, zero, AND_A17_B0);

    wire AND_A18_B0;
    and and_a18_b0(AND_A18_B0, A[18], B[0]);
    wire P_A18_B0, Cout_A18_B0;
    half_adder add_a18_b0(P_A18_B0, Cout_A18_B0, zero, AND_A18_B0);

    wire AND_A19_B0;
    and and_a19_b0(AND_A19_B0, A[19], B[0]);
    wire P_A19_B0, Cout_A19_B0;
    half_adder add_a19_b0(P_A19_B0, Cout_A19_B0, zero, AND_A19_B0);

    wire AND_A20_B0;
    and and_a20_b0(AND_A20_B0, A[20], B[0]);
    wire P_A20_B0, Cout_A20_B0;
    half_adder add_a20_b0(P_A20_B0, Cout_A20_B0, zero, AND_A20_B0);

    wire AND_A21_B0;
    and and_a21_b0(AND_A21_B0, A[21], B[0]);
    wire P_A21_B0, Cout_A21_B0;
    half_adder add_a21_b0(P_A21_B0, Cout_A21_B0, zero, AND_A21_B0);

    wire AND_A22_B0;
    and and_a22_b0(AND_A22_B0, A[22], B[0]);
    wire P_A22_B0, Cout_A22_B0;
    half_adder add_a22_b0(P_A22_B0, Cout_A22_B0, zero, AND_A22_B0);

    wire AND_A23_B0;
    and and_a23_b0(AND_A23_B0, A[23], B[0]);
    wire P_A23_B0, Cout_A23_B0;
    half_adder add_a23_b0(P_A23_B0, Cout_A23_B0, zero, AND_A23_B0);

    wire AND_A24_B0;
    and and_a24_b0(AND_A24_B0, A[24], B[0]);
    wire P_A24_B0, Cout_A24_B0;
    half_adder add_a24_b0(P_A24_B0, Cout_A24_B0, zero, AND_A24_B0);

    wire AND_A25_B0;
    and and_a25_b0(AND_A25_B0, A[25], B[0]);
    wire P_A25_B0, Cout_A25_B0;
    half_adder add_a25_b0(P_A25_B0, Cout_A25_B0, zero, AND_A25_B0);

    wire AND_A26_B0;
    and and_a26_b0(AND_A26_B0, A[26], B[0]);
    wire P_A26_B0, Cout_A26_B0;
    half_adder add_a26_b0(P_A26_B0, Cout_A26_B0, zero, AND_A26_B0);

    wire AND_A27_B0;
    and and_a27_b0(AND_A27_B0, A[27], B[0]);
    wire P_A27_B0, Cout_A27_B0;
    half_adder add_a27_b0(P_A27_B0, Cout_A27_B0, zero, AND_A27_B0);

    wire AND_A28_B0;
    and and_a28_b0(AND_A28_B0, A[28], B[0]);
    wire P_A28_B0, Cout_A28_B0;
    half_adder add_a28_b0(P_A28_B0, Cout_A28_B0, zero, AND_A28_B0);

    wire AND_A29_B0;
    and and_a29_b0(AND_A29_B0, A[29], B[0]);
    wire P_A29_B0, Cout_A29_B0;
    half_adder add_a29_b0(P_A29_B0, Cout_A29_B0, zero, AND_A29_B0);

    wire AND_A30_B0;
    and and_a30_b0(AND_A30_B0, A[30], B[0]);
    wire P_A30_B0, Cout_A30_B0;
    half_adder add_a30_b0(P_A30_B0, Cout_A30_B0, zero, AND_A30_B0);

    wire AND_A31_B0;
    nand and_a31_b0(AND_A31_B0, A[31], B[0]);
    wire P_A31_B0, Cout_A31_B0;
    half_adder add_a31_b0(P_A31_B0, Cout_A31_B0, zero, AND_A31_B0);

    wire AND_A0_B1;
    and and_a0_b1(AND_A0_B1, A[0], B[1]);
    wire P_A0_B1, Cout_A0_B1;
    full_adder add_a0_b1(P_A0_B1, Cout_A0_B1, P_A1_B0, AND_A0_B1, Cout_A0_B0);

    wire AND_A1_B1;
    and and_a1_b1(AND_A1_B1, A[1], B[1]);
    wire P_A1_B1, Cout_A1_B1;
    full_adder add_a1_b1(P_A1_B1, Cout_A1_B1, P_A2_B0, AND_A1_B1, Cout_A1_B0);

    wire AND_A2_B1;
    and and_a2_b1(AND_A2_B1, A[2], B[1]);
    wire P_A2_B1, Cout_A2_B1;
    full_adder add_a2_b1(P_A2_B1, Cout_A2_B1, P_A3_B0, AND_A2_B1, Cout_A2_B0);

    wire AND_A3_B1;
    and and_a3_b1(AND_A3_B1, A[3], B[1]);
    wire P_A3_B1, Cout_A3_B1;
    full_adder add_a3_b1(P_A3_B1, Cout_A3_B1, P_A4_B0, AND_A3_B1, Cout_A3_B0);

    wire AND_A4_B1;
    and and_a4_b1(AND_A4_B1, A[4], B[1]);
    wire P_A4_B1, Cout_A4_B1;
    full_adder add_a4_b1(P_A4_B1, Cout_A4_B1, P_A5_B0, AND_A4_B1, Cout_A4_B0);

    wire AND_A5_B1;
    and and_a5_b1(AND_A5_B1, A[5], B[1]);
    wire P_A5_B1, Cout_A5_B1;
    full_adder add_a5_b1(P_A5_B1, Cout_A5_B1, P_A6_B0, AND_A5_B1, Cout_A5_B0);

    wire AND_A6_B1;
    and and_a6_b1(AND_A6_B1, A[6], B[1]);
    wire P_A6_B1, Cout_A6_B1;
    full_adder add_a6_b1(P_A6_B1, Cout_A6_B1, P_A7_B0, AND_A6_B1, Cout_A6_B0);

    wire AND_A7_B1;
    and and_a7_b1(AND_A7_B1, A[7], B[1]);
    wire P_A7_B1, Cout_A7_B1;
    full_adder add_a7_b1(P_A7_B1, Cout_A7_B1, P_A8_B0, AND_A7_B1, Cout_A7_B0);

    wire AND_A8_B1;
    and and_a8_b1(AND_A8_B1, A[8], B[1]);
    wire P_A8_B1, Cout_A8_B1;
    full_adder add_a8_b1(P_A8_B1, Cout_A8_B1, P_A9_B0, AND_A8_B1, Cout_A8_B0);

    wire AND_A9_B1;
    and and_a9_b1(AND_A9_B1, A[9], B[1]);
    wire P_A9_B1, Cout_A9_B1;
    full_adder add_a9_b1(P_A9_B1, Cout_A9_B1, P_A10_B0, AND_A9_B1, Cout_A9_B0);

    wire AND_A10_B1;
    and and_a10_b1(AND_A10_B1, A[10], B[1]);
    wire P_A10_B1, Cout_A10_B1;
    full_adder add_a10_b1(P_A10_B1, Cout_A10_B1, P_A11_B0, AND_A10_B1, Cout_A10_B0);

    wire AND_A11_B1;
    and and_a11_b1(AND_A11_B1, A[11], B[1]);
    wire P_A11_B1, Cout_A11_B1;
    full_adder add_a11_b1(P_A11_B1, Cout_A11_B1, P_A12_B0, AND_A11_B1, Cout_A11_B0);

    wire AND_A12_B1;
    and and_a12_b1(AND_A12_B1, A[12], B[1]);
    wire P_A12_B1, Cout_A12_B1;
    full_adder add_a12_b1(P_A12_B1, Cout_A12_B1, P_A13_B0, AND_A12_B1, Cout_A12_B0);

    wire AND_A13_B1;
    and and_a13_b1(AND_A13_B1, A[13], B[1]);
    wire P_A13_B1, Cout_A13_B1;
    full_adder add_a13_b1(P_A13_B1, Cout_A13_B1, P_A14_B0, AND_A13_B1, Cout_A13_B0);

    wire AND_A14_B1;
    and and_a14_b1(AND_A14_B1, A[14], B[1]);
    wire P_A14_B1, Cout_A14_B1;
    full_adder add_a14_b1(P_A14_B1, Cout_A14_B1, P_A15_B0, AND_A14_B1, Cout_A14_B0);

    wire AND_A15_B1;
    and and_a15_b1(AND_A15_B1, A[15], B[1]);
    wire P_A15_B1, Cout_A15_B1;
    full_adder add_a15_b1(P_A15_B1, Cout_A15_B1, P_A16_B0, AND_A15_B1, Cout_A15_B0);

    wire AND_A16_B1;
    and and_a16_b1(AND_A16_B1, A[16], B[1]);
    wire P_A16_B1, Cout_A16_B1;
    full_adder add_a16_b1(P_A16_B1, Cout_A16_B1, P_A17_B0, AND_A16_B1, Cout_A16_B0);

    wire AND_A17_B1;
    and and_a17_b1(AND_A17_B1, A[17], B[1]);
    wire P_A17_B1, Cout_A17_B1;
    full_adder add_a17_b1(P_A17_B1, Cout_A17_B1, P_A18_B0, AND_A17_B1, Cout_A17_B0);

    wire AND_A18_B1;
    and and_a18_b1(AND_A18_B1, A[18], B[1]);
    wire P_A18_B1, Cout_A18_B1;
    full_adder add_a18_b1(P_A18_B1, Cout_A18_B1, P_A19_B0, AND_A18_B1, Cout_A18_B0);

    wire AND_A19_B1;
    and and_a19_b1(AND_A19_B1, A[19], B[1]);
    wire P_A19_B1, Cout_A19_B1;
    full_adder add_a19_b1(P_A19_B1, Cout_A19_B1, P_A20_B0, AND_A19_B1, Cout_A19_B0);

    wire AND_A20_B1;
    and and_a20_b1(AND_A20_B1, A[20], B[1]);
    wire P_A20_B1, Cout_A20_B1;
    full_adder add_a20_b1(P_A20_B1, Cout_A20_B1, P_A21_B0, AND_A20_B1, Cout_A20_B0);

    wire AND_A21_B1;
    and and_a21_b1(AND_A21_B1, A[21], B[1]);
    wire P_A21_B1, Cout_A21_B1;
    full_adder add_a21_b1(P_A21_B1, Cout_A21_B1, P_A22_B0, AND_A21_B1, Cout_A21_B0);

    wire AND_A22_B1;
    and and_a22_b1(AND_A22_B1, A[22], B[1]);
    wire P_A22_B1, Cout_A22_B1;
    full_adder add_a22_b1(P_A22_B1, Cout_A22_B1, P_A23_B0, AND_A22_B1, Cout_A22_B0);

    wire AND_A23_B1;
    and and_a23_b1(AND_A23_B1, A[23], B[1]);
    wire P_A23_B1, Cout_A23_B1;
    full_adder add_a23_b1(P_A23_B1, Cout_A23_B1, P_A24_B0, AND_A23_B1, Cout_A23_B0);

    wire AND_A24_B1;
    and and_a24_b1(AND_A24_B1, A[24], B[1]);
    wire P_A24_B1, Cout_A24_B1;
    full_adder add_a24_b1(P_A24_B1, Cout_A24_B1, P_A25_B0, AND_A24_B1, Cout_A24_B0);

    wire AND_A25_B1;
    and and_a25_b1(AND_A25_B1, A[25], B[1]);
    wire P_A25_B1, Cout_A25_B1;
    full_adder add_a25_b1(P_A25_B1, Cout_A25_B1, P_A26_B0, AND_A25_B1, Cout_A25_B0);

    wire AND_A26_B1;
    and and_a26_b1(AND_A26_B1, A[26], B[1]);
    wire P_A26_B1, Cout_A26_B1;
    full_adder add_a26_b1(P_A26_B1, Cout_A26_B1, P_A27_B0, AND_A26_B1, Cout_A26_B0);

    wire AND_A27_B1;
    and and_a27_b1(AND_A27_B1, A[27], B[1]);
    wire P_A27_B1, Cout_A27_B1;
    full_adder add_a27_b1(P_A27_B1, Cout_A27_B1, P_A28_B0, AND_A27_B1, Cout_A27_B0);

    wire AND_A28_B1;
    and and_a28_b1(AND_A28_B1, A[28], B[1]);
    wire P_A28_B1, Cout_A28_B1;
    full_adder add_a28_b1(P_A28_B1, Cout_A28_B1, P_A29_B0, AND_A28_B1, Cout_A28_B0);

    wire AND_A29_B1;
    and and_a29_b1(AND_A29_B1, A[29], B[1]);
    wire P_A29_B1, Cout_A29_B1;
    full_adder add_a29_b1(P_A29_B1, Cout_A29_B1, P_A30_B0, AND_A29_B1, Cout_A29_B0);

    wire AND_A30_B1;
    and and_a30_b1(AND_A30_B1, A[30], B[1]);
    wire P_A30_B1, Cout_A30_B1;
    full_adder add_a30_b1(P_A30_B1, Cout_A30_B1, P_A31_B0, AND_A30_B1, Cout_A30_B0);

    wire AND_A31_B1;
    nand and_a31_b1(AND_A31_B1, A[31], B[1]);
    wire P_A31_B1, Cout_A31_B1;
    wire single_one;
    assign single_one = 1'b1;
    full_adder add_a31_b1(P_A31_B1, Cout_A31_B1, AND_A31_B1, Cout_A31_B0, single_one);

    wire AND_A0_B2;
    and and_a0_b2(AND_A0_B2, A[0], B[2]);
    wire P_A0_B2, Cout_A0_B2;
    full_adder add_a0_b2(P_A0_B2, Cout_A0_B2, P_A1_B1, AND_A0_B2, Cout_A0_B1);

    wire AND_A1_B2;
    and and_a1_b2(AND_A1_B2, A[1], B[2]);
    wire P_A1_B2, Cout_A1_B2;
    full_adder add_a1_b2(P_A1_B2, Cout_A1_B2, P_A2_B1, AND_A1_B2, Cout_A1_B1);

    wire AND_A2_B2;
    and and_a2_b2(AND_A2_B2, A[2], B[2]);
    wire P_A2_B2, Cout_A2_B2;
    full_adder add_a2_b2(P_A2_B2, Cout_A2_B2, P_A3_B1, AND_A2_B2, Cout_A2_B1);

    wire AND_A3_B2;
    and and_a3_b2(AND_A3_B2, A[3], B[2]);
    wire P_A3_B2, Cout_A3_B2;
    full_adder add_a3_b2(P_A3_B2, Cout_A3_B2, P_A4_B1, AND_A3_B2, Cout_A3_B1);

    wire AND_A4_B2;
    and and_a4_b2(AND_A4_B2, A[4], B[2]);
    wire P_A4_B2, Cout_A4_B2;
    full_adder add_a4_b2(P_A4_B2, Cout_A4_B2, P_A5_B1, AND_A4_B2, Cout_A4_B1);

    wire AND_A5_B2;
    and and_a5_b2(AND_A5_B2, A[5], B[2]);
    wire P_A5_B2, Cout_A5_B2;
    full_adder add_a5_b2(P_A5_B2, Cout_A5_B2, P_A6_B1, AND_A5_B2, Cout_A5_B1);

    wire AND_A6_B2;
    and and_a6_b2(AND_A6_B2, A[6], B[2]);
    wire P_A6_B2, Cout_A6_B2;
    full_adder add_a6_b2(P_A6_B2, Cout_A6_B2, P_A7_B1, AND_A6_B2, Cout_A6_B1);

    wire AND_A7_B2;
    and and_a7_b2(AND_A7_B2, A[7], B[2]);
    wire P_A7_B2, Cout_A7_B2;
    full_adder add_a7_b2(P_A7_B2, Cout_A7_B2, P_A8_B1, AND_A7_B2, Cout_A7_B1);

    wire AND_A8_B2;
    and and_a8_b2(AND_A8_B2, A[8], B[2]);
    wire P_A8_B2, Cout_A8_B2;
    full_adder add_a8_b2(P_A8_B2, Cout_A8_B2, P_A9_B1, AND_A8_B2, Cout_A8_B1);

    wire AND_A9_B2;
    and and_a9_b2(AND_A9_B2, A[9], B[2]);
    wire P_A9_B2, Cout_A9_B2;
    full_adder add_a9_b2(P_A9_B2, Cout_A9_B2, P_A10_B1, AND_A9_B2, Cout_A9_B1);

    wire AND_A10_B2;
    and and_a10_b2(AND_A10_B2, A[10], B[2]);
    wire P_A10_B2, Cout_A10_B2;
    full_adder add_a10_b2(P_A10_B2, Cout_A10_B2, P_A11_B1, AND_A10_B2, Cout_A10_B1);

    wire AND_A11_B2;
    and and_a11_b2(AND_A11_B2, A[11], B[2]);
    wire P_A11_B2, Cout_A11_B2;
    full_adder add_a11_b2(P_A11_B2, Cout_A11_B2, P_A12_B1, AND_A11_B2, Cout_A11_B1);

    wire AND_A12_B2;
    and and_a12_b2(AND_A12_B2, A[12], B[2]);
    wire P_A12_B2, Cout_A12_B2;
    full_adder add_a12_b2(P_A12_B2, Cout_A12_B2, P_A13_B1, AND_A12_B2, Cout_A12_B1);

    wire AND_A13_B2;
    and and_a13_b2(AND_A13_B2, A[13], B[2]);
    wire P_A13_B2, Cout_A13_B2;
    full_adder add_a13_b2(P_A13_B2, Cout_A13_B2, P_A14_B1, AND_A13_B2, Cout_A13_B1);

    wire AND_A14_B2;
    and and_a14_b2(AND_A14_B2, A[14], B[2]);
    wire P_A14_B2, Cout_A14_B2;
    full_adder add_a14_b2(P_A14_B2, Cout_A14_B2, P_A15_B1, AND_A14_B2, Cout_A14_B1);

    wire AND_A15_B2;
    and and_a15_b2(AND_A15_B2, A[15], B[2]);
    wire P_A15_B2, Cout_A15_B2;
    full_adder add_a15_b2(P_A15_B2, Cout_A15_B2, P_A16_B1, AND_A15_B2, Cout_A15_B1);

    wire AND_A16_B2;
    and and_a16_b2(AND_A16_B2, A[16], B[2]);
    wire P_A16_B2, Cout_A16_B2;
    full_adder add_a16_b2(P_A16_B2, Cout_A16_B2, P_A17_B1, AND_A16_B2, Cout_A16_B1);

    wire AND_A17_B2;
    and and_a17_b2(AND_A17_B2, A[17], B[2]);
    wire P_A17_B2, Cout_A17_B2;
    full_adder add_a17_b2(P_A17_B2, Cout_A17_B2, P_A18_B1, AND_A17_B2, Cout_A17_B1);

    wire AND_A18_B2;
    and and_a18_b2(AND_A18_B2, A[18], B[2]);
    wire P_A18_B2, Cout_A18_B2;
    full_adder add_a18_b2(P_A18_B2, Cout_A18_B2, P_A19_B1, AND_A18_B2, Cout_A18_B1);

    wire AND_A19_B2;
    and and_a19_b2(AND_A19_B2, A[19], B[2]);
    wire P_A19_B2, Cout_A19_B2;
    full_adder add_a19_b2(P_A19_B2, Cout_A19_B2, P_A20_B1, AND_A19_B2, Cout_A19_B1);

    wire AND_A20_B2;
    and and_a20_b2(AND_A20_B2, A[20], B[2]);
    wire P_A20_B2, Cout_A20_B2;
    full_adder add_a20_b2(P_A20_B2, Cout_A20_B2, P_A21_B1, AND_A20_B2, Cout_A20_B1);

    wire AND_A21_B2;
    and and_a21_b2(AND_A21_B2, A[21], B[2]);
    wire P_A21_B2, Cout_A21_B2;
    full_adder add_a21_b2(P_A21_B2, Cout_A21_B2, P_A22_B1, AND_A21_B2, Cout_A21_B1);

    wire AND_A22_B2;
    and and_a22_b2(AND_A22_B2, A[22], B[2]);
    wire P_A22_B2, Cout_A22_B2;
    full_adder add_a22_b2(P_A22_B2, Cout_A22_B2, P_A23_B1, AND_A22_B2, Cout_A22_B1);

    wire AND_A23_B2;
    and and_a23_b2(AND_A23_B2, A[23], B[2]);
    wire P_A23_B2, Cout_A23_B2;
    full_adder add_a23_b2(P_A23_B2, Cout_A23_B2, P_A24_B1, AND_A23_B2, Cout_A23_B1);

    wire AND_A24_B2;
    and and_a24_b2(AND_A24_B2, A[24], B[2]);
    wire P_A24_B2, Cout_A24_B2;
    full_adder add_a24_b2(P_A24_B2, Cout_A24_B2, P_A25_B1, AND_A24_B2, Cout_A24_B1);

    wire AND_A25_B2;
    and and_a25_b2(AND_A25_B2, A[25], B[2]);
    wire P_A25_B2, Cout_A25_B2;
    full_adder add_a25_b2(P_A25_B2, Cout_A25_B2, P_A26_B1, AND_A25_B2, Cout_A25_B1);

    wire AND_A26_B2;
    and and_a26_b2(AND_A26_B2, A[26], B[2]);
    wire P_A26_B2, Cout_A26_B2;
    full_adder add_a26_b2(P_A26_B2, Cout_A26_B2, P_A27_B1, AND_A26_B2, Cout_A26_B1);

    wire AND_A27_B2;
    and and_a27_b2(AND_A27_B2, A[27], B[2]);
    wire P_A27_B2, Cout_A27_B2;
    full_adder add_a27_b2(P_A27_B2, Cout_A27_B2, P_A28_B1, AND_A27_B2, Cout_A27_B1);

    wire AND_A28_B2;
    and and_a28_b2(AND_A28_B2, A[28], B[2]);
    wire P_A28_B2, Cout_A28_B2;
    full_adder add_a28_b2(P_A28_B2, Cout_A28_B2, P_A29_B1, AND_A28_B2, Cout_A28_B1);

    wire AND_A29_B2;
    and and_a29_b2(AND_A29_B2, A[29], B[2]);
    wire P_A29_B2, Cout_A29_B2;
    full_adder add_a29_b2(P_A29_B2, Cout_A29_B2, P_A30_B1, AND_A29_B2, Cout_A29_B1);

    wire AND_A30_B2;
    and and_a30_b2(AND_A30_B2, A[30], B[2]);
    wire P_A30_B2, Cout_A30_B2;
    full_adder add_a30_b2(P_A30_B2, Cout_A30_B2, P_A31_B1, AND_A30_B2, Cout_A30_B1);

    wire AND_A31_B2;
    nand and_a31_b2(AND_A31_B2, A[31], B[2]);
    wire P_A31_B2, Cout_A31_B2;
    half_adder add_a31_b2(P_A31_B2, Cout_A31_B2, AND_A31_B2, Cout_A31_B1);

    wire AND_A0_B3;
    and and_a0_b3(AND_A0_B3, A[0], B[3]);
    wire P_A0_B3, Cout_A0_B3;
    full_adder add_a0_b3(P_A0_B3, Cout_A0_B3, P_A1_B2, AND_A0_B3, Cout_A0_B2);

    wire AND_A1_B3;
    and and_a1_b3(AND_A1_B3, A[1], B[3]);
    wire P_A1_B3, Cout_A1_B3;
    full_adder add_a1_b3(P_A1_B3, Cout_A1_B3, P_A2_B2, AND_A1_B3, Cout_A1_B2);

    wire AND_A2_B3;
    and and_a2_b3(AND_A2_B3, A[2], B[3]);
    wire P_A2_B3, Cout_A2_B3;
    full_adder add_a2_b3(P_A2_B3, Cout_A2_B3, P_A3_B2, AND_A2_B3, Cout_A2_B2);

    wire AND_A3_B3;
    and and_a3_b3(AND_A3_B3, A[3], B[3]);
    wire P_A3_B3, Cout_A3_B3;
    full_adder add_a3_b3(P_A3_B3, Cout_A3_B3, P_A4_B2, AND_A3_B3, Cout_A3_B2);

    wire AND_A4_B3;
    and and_a4_b3(AND_A4_B3, A[4], B[3]);
    wire P_A4_B3, Cout_A4_B3;
    full_adder add_a4_b3(P_A4_B3, Cout_A4_B3, P_A5_B2, AND_A4_B3, Cout_A4_B2);

    wire AND_A5_B3;
    and and_a5_b3(AND_A5_B3, A[5], B[3]);
    wire P_A5_B3, Cout_A5_B3;
    full_adder add_a5_b3(P_A5_B3, Cout_A5_B3, P_A6_B2, AND_A5_B3, Cout_A5_B2);

    wire AND_A6_B3;
    and and_a6_b3(AND_A6_B3, A[6], B[3]);
    wire P_A6_B3, Cout_A6_B3;
    full_adder add_a6_b3(P_A6_B3, Cout_A6_B3, P_A7_B2, AND_A6_B3, Cout_A6_B2);

    wire AND_A7_B3;
    and and_a7_b3(AND_A7_B3, A[7], B[3]);
    wire P_A7_B3, Cout_A7_B3;
    full_adder add_a7_b3(P_A7_B3, Cout_A7_B3, P_A8_B2, AND_A7_B3, Cout_A7_B2);

    wire AND_A8_B3;
    and and_a8_b3(AND_A8_B3, A[8], B[3]);
    wire P_A8_B3, Cout_A8_B3;
    full_adder add_a8_b3(P_A8_B3, Cout_A8_B3, P_A9_B2, AND_A8_B3, Cout_A8_B2);

    wire AND_A9_B3;
    and and_a9_b3(AND_A9_B3, A[9], B[3]);
    wire P_A9_B3, Cout_A9_B3;
    full_adder add_a9_b3(P_A9_B3, Cout_A9_B3, P_A10_B2, AND_A9_B3, Cout_A9_B2);

    wire AND_A10_B3;
    and and_a10_b3(AND_A10_B3, A[10], B[3]);
    wire P_A10_B3, Cout_A10_B3;
    full_adder add_a10_b3(P_A10_B3, Cout_A10_B3, P_A11_B2, AND_A10_B3, Cout_A10_B2);

    wire AND_A11_B3;
    and and_a11_b3(AND_A11_B3, A[11], B[3]);
    wire P_A11_B3, Cout_A11_B3;
    full_adder add_a11_b3(P_A11_B3, Cout_A11_B3, P_A12_B2, AND_A11_B3, Cout_A11_B2);

    wire AND_A12_B3;
    and and_a12_b3(AND_A12_B3, A[12], B[3]);
    wire P_A12_B3, Cout_A12_B3;
    full_adder add_a12_b3(P_A12_B3, Cout_A12_B3, P_A13_B2, AND_A12_B3, Cout_A12_B2);

    wire AND_A13_B3;
    and and_a13_b3(AND_A13_B3, A[13], B[3]);
    wire P_A13_B3, Cout_A13_B3;
    full_adder add_a13_b3(P_A13_B3, Cout_A13_B3, P_A14_B2, AND_A13_B3, Cout_A13_B2);

    wire AND_A14_B3;
    and and_a14_b3(AND_A14_B3, A[14], B[3]);
    wire P_A14_B3, Cout_A14_B3;
    full_adder add_a14_b3(P_A14_B3, Cout_A14_B3, P_A15_B2, AND_A14_B3, Cout_A14_B2);

    wire AND_A15_B3;
    and and_a15_b3(AND_A15_B3, A[15], B[3]);
    wire P_A15_B3, Cout_A15_B3;
    full_adder add_a15_b3(P_A15_B3, Cout_A15_B3, P_A16_B2, AND_A15_B3, Cout_A15_B2);

    wire AND_A16_B3;
    and and_a16_b3(AND_A16_B3, A[16], B[3]);
    wire P_A16_B3, Cout_A16_B3;
    full_adder add_a16_b3(P_A16_B3, Cout_A16_B3, P_A17_B2, AND_A16_B3, Cout_A16_B2);

    wire AND_A17_B3;
    and and_a17_b3(AND_A17_B3, A[17], B[3]);
    wire P_A17_B3, Cout_A17_B3;
    full_adder add_a17_b3(P_A17_B3, Cout_A17_B3, P_A18_B2, AND_A17_B3, Cout_A17_B2);

    wire AND_A18_B3;
    and and_a18_b3(AND_A18_B3, A[18], B[3]);
    wire P_A18_B3, Cout_A18_B3;
    full_adder add_a18_b3(P_A18_B3, Cout_A18_B3, P_A19_B2, AND_A18_B3, Cout_A18_B2);

    wire AND_A19_B3;
    and and_a19_b3(AND_A19_B3, A[19], B[3]);
    wire P_A19_B3, Cout_A19_B3;
    full_adder add_a19_b3(P_A19_B3, Cout_A19_B3, P_A20_B2, AND_A19_B3, Cout_A19_B2);

    wire AND_A20_B3;
    and and_a20_b3(AND_A20_B3, A[20], B[3]);
    wire P_A20_B3, Cout_A20_B3;
    full_adder add_a20_b3(P_A20_B3, Cout_A20_B3, P_A21_B2, AND_A20_B3, Cout_A20_B2);

    wire AND_A21_B3;
    and and_a21_b3(AND_A21_B3, A[21], B[3]);
    wire P_A21_B3, Cout_A21_B3;
    full_adder add_a21_b3(P_A21_B3, Cout_A21_B3, P_A22_B2, AND_A21_B3, Cout_A21_B2);

    wire AND_A22_B3;
    and and_a22_b3(AND_A22_B3, A[22], B[3]);
    wire P_A22_B3, Cout_A22_B3;
    full_adder add_a22_b3(P_A22_B3, Cout_A22_B3, P_A23_B2, AND_A22_B3, Cout_A22_B2);

    wire AND_A23_B3;
    and and_a23_b3(AND_A23_B3, A[23], B[3]);
    wire P_A23_B3, Cout_A23_B3;
    full_adder add_a23_b3(P_A23_B3, Cout_A23_B3, P_A24_B2, AND_A23_B3, Cout_A23_B2);

    wire AND_A24_B3;
    and and_a24_b3(AND_A24_B3, A[24], B[3]);
    wire P_A24_B3, Cout_A24_B3;
    full_adder add_a24_b3(P_A24_B3, Cout_A24_B3, P_A25_B2, AND_A24_B3, Cout_A24_B2);

    wire AND_A25_B3;
    and and_a25_b3(AND_A25_B3, A[25], B[3]);
    wire P_A25_B3, Cout_A25_B3;
    full_adder add_a25_b3(P_A25_B3, Cout_A25_B3, P_A26_B2, AND_A25_B3, Cout_A25_B2);

    wire AND_A26_B3;
    and and_a26_b3(AND_A26_B3, A[26], B[3]);
    wire P_A26_B3, Cout_A26_B3;
    full_adder add_a26_b3(P_A26_B3, Cout_A26_B3, P_A27_B2, AND_A26_B3, Cout_A26_B2);

    wire AND_A27_B3;
    and and_a27_b3(AND_A27_B3, A[27], B[3]);
    wire P_A27_B3, Cout_A27_B3;
    full_adder add_a27_b3(P_A27_B3, Cout_A27_B3, P_A28_B2, AND_A27_B3, Cout_A27_B2);

    wire AND_A28_B3;
    and and_a28_b3(AND_A28_B3, A[28], B[3]);
    wire P_A28_B3, Cout_A28_B3;
    full_adder add_a28_b3(P_A28_B3, Cout_A28_B3, P_A29_B2, AND_A28_B3, Cout_A28_B2);

    wire AND_A29_B3;
    and and_a29_b3(AND_A29_B3, A[29], B[3]);
    wire P_A29_B3, Cout_A29_B3;
    full_adder add_a29_b3(P_A29_B3, Cout_A29_B3, P_A30_B2, AND_A29_B3, Cout_A29_B2);

    wire AND_A30_B3;
    and and_a30_b3(AND_A30_B3, A[30], B[3]);
    wire P_A30_B3, Cout_A30_B3;
    full_adder add_a30_b3(P_A30_B3, Cout_A30_B3, P_A31_B2, AND_A30_B3, Cout_A30_B2);

    wire AND_A31_B3;
    nand and_a31_b3(AND_A31_B3, A[31], B[3]);
    wire P_A31_B3, Cout_A31_B3;
    half_adder add_a31_b3(P_A31_B3, Cout_A31_B3, AND_A31_B3, Cout_A31_B2);

    wire AND_A0_B4;
    and and_a0_b4(AND_A0_B4, A[0], B[4]);
    wire P_A0_B4, Cout_A0_B4;
    full_adder add_a0_b4(P_A0_B4, Cout_A0_B4, P_A1_B3, AND_A0_B4, Cout_A0_B3);

    wire AND_A1_B4;
    and and_a1_b4(AND_A1_B4, A[1], B[4]);
    wire P_A1_B4, Cout_A1_B4;
    full_adder add_a1_b4(P_A1_B4, Cout_A1_B4, P_A2_B3, AND_A1_B4, Cout_A1_B3);

    wire AND_A2_B4;
    and and_a2_b4(AND_A2_B4, A[2], B[4]);
    wire P_A2_B4, Cout_A2_B4;
    full_adder add_a2_b4(P_A2_B4, Cout_A2_B4, P_A3_B3, AND_A2_B4, Cout_A2_B3);

    wire AND_A3_B4;
    and and_a3_b4(AND_A3_B4, A[3], B[4]);
    wire P_A3_B4, Cout_A3_B4;
    full_adder add_a3_b4(P_A3_B4, Cout_A3_B4, P_A4_B3, AND_A3_B4, Cout_A3_B3);

    wire AND_A4_B4;
    and and_a4_b4(AND_A4_B4, A[4], B[4]);
    wire P_A4_B4, Cout_A4_B4;
    full_adder add_a4_b4(P_A4_B4, Cout_A4_B4, P_A5_B3, AND_A4_B4, Cout_A4_B3);

    wire AND_A5_B4;
    and and_a5_b4(AND_A5_B4, A[5], B[4]);
    wire P_A5_B4, Cout_A5_B4;
    full_adder add_a5_b4(P_A5_B4, Cout_A5_B4, P_A6_B3, AND_A5_B4, Cout_A5_B3);

    wire AND_A6_B4;
    and and_a6_b4(AND_A6_B4, A[6], B[4]);
    wire P_A6_B4, Cout_A6_B4;
    full_adder add_a6_b4(P_A6_B4, Cout_A6_B4, P_A7_B3, AND_A6_B4, Cout_A6_B3);

    wire AND_A7_B4;
    and and_a7_b4(AND_A7_B4, A[7], B[4]);
    wire P_A7_B4, Cout_A7_B4;
    full_adder add_a7_b4(P_A7_B4, Cout_A7_B4, P_A8_B3, AND_A7_B4, Cout_A7_B3);

    wire AND_A8_B4;
    and and_a8_b4(AND_A8_B4, A[8], B[4]);
    wire P_A8_B4, Cout_A8_B4;
    full_adder add_a8_b4(P_A8_B4, Cout_A8_B4, P_A9_B3, AND_A8_B4, Cout_A8_B3);

    wire AND_A9_B4;
    and and_a9_b4(AND_A9_B4, A[9], B[4]);
    wire P_A9_B4, Cout_A9_B4;
    full_adder add_a9_b4(P_A9_B4, Cout_A9_B4, P_A10_B3, AND_A9_B4, Cout_A9_B3);

    wire AND_A10_B4;
    and and_a10_b4(AND_A10_B4, A[10], B[4]);
    wire P_A10_B4, Cout_A10_B4;
    full_adder add_a10_b4(P_A10_B4, Cout_A10_B4, P_A11_B3, AND_A10_B4, Cout_A10_B3);

    wire AND_A11_B4;
    and and_a11_b4(AND_A11_B4, A[11], B[4]);
    wire P_A11_B4, Cout_A11_B4;
    full_adder add_a11_b4(P_A11_B4, Cout_A11_B4, P_A12_B3, AND_A11_B4, Cout_A11_B3);

    wire AND_A12_B4;
    and and_a12_b4(AND_A12_B4, A[12], B[4]);
    wire P_A12_B4, Cout_A12_B4;
    full_adder add_a12_b4(P_A12_B4, Cout_A12_B4, P_A13_B3, AND_A12_B4, Cout_A12_B3);

    wire AND_A13_B4;
    and and_a13_b4(AND_A13_B4, A[13], B[4]);
    wire P_A13_B4, Cout_A13_B4;
    full_adder add_a13_b4(P_A13_B4, Cout_A13_B4, P_A14_B3, AND_A13_B4, Cout_A13_B3);

    wire AND_A14_B4;
    and and_a14_b4(AND_A14_B4, A[14], B[4]);
    wire P_A14_B4, Cout_A14_B4;
    full_adder add_a14_b4(P_A14_B4, Cout_A14_B4, P_A15_B3, AND_A14_B4, Cout_A14_B3);

    wire AND_A15_B4;
    and and_a15_b4(AND_A15_B4, A[15], B[4]);
    wire P_A15_B4, Cout_A15_B4;
    full_adder add_a15_b4(P_A15_B4, Cout_A15_B4, P_A16_B3, AND_A15_B4, Cout_A15_B3);

    wire AND_A16_B4;
    and and_a16_b4(AND_A16_B4, A[16], B[4]);
    wire P_A16_B4, Cout_A16_B4;
    full_adder add_a16_b4(P_A16_B4, Cout_A16_B4, P_A17_B3, AND_A16_B4, Cout_A16_B3);

    wire AND_A17_B4;
    and and_a17_b4(AND_A17_B4, A[17], B[4]);
    wire P_A17_B4, Cout_A17_B4;
    full_adder add_a17_b4(P_A17_B4, Cout_A17_B4, P_A18_B3, AND_A17_B4, Cout_A17_B3);

    wire AND_A18_B4;
    and and_a18_b4(AND_A18_B4, A[18], B[4]);
    wire P_A18_B4, Cout_A18_B4;
    full_adder add_a18_b4(P_A18_B4, Cout_A18_B4, P_A19_B3, AND_A18_B4, Cout_A18_B3);

    wire AND_A19_B4;
    and and_a19_b4(AND_A19_B4, A[19], B[4]);
    wire P_A19_B4, Cout_A19_B4;
    full_adder add_a19_b4(P_A19_B4, Cout_A19_B4, P_A20_B3, AND_A19_B4, Cout_A19_B3);

    wire AND_A20_B4;
    and and_a20_b4(AND_A20_B4, A[20], B[4]);
    wire P_A20_B4, Cout_A20_B4;
    full_adder add_a20_b4(P_A20_B4, Cout_A20_B4, P_A21_B3, AND_A20_B4, Cout_A20_B3);

    wire AND_A21_B4;
    and and_a21_b4(AND_A21_B4, A[21], B[4]);
    wire P_A21_B4, Cout_A21_B4;
    full_adder add_a21_b4(P_A21_B4, Cout_A21_B4, P_A22_B3, AND_A21_B4, Cout_A21_B3);

    wire AND_A22_B4;
    and and_a22_b4(AND_A22_B4, A[22], B[4]);
    wire P_A22_B4, Cout_A22_B4;
    full_adder add_a22_b4(P_A22_B4, Cout_A22_B4, P_A23_B3, AND_A22_B4, Cout_A22_B3);

    wire AND_A23_B4;
    and and_a23_b4(AND_A23_B4, A[23], B[4]);
    wire P_A23_B4, Cout_A23_B4;
    full_adder add_a23_b4(P_A23_B4, Cout_A23_B4, P_A24_B3, AND_A23_B4, Cout_A23_B3);

    wire AND_A24_B4;
    and and_a24_b4(AND_A24_B4, A[24], B[4]);
    wire P_A24_B4, Cout_A24_B4;
    full_adder add_a24_b4(P_A24_B4, Cout_A24_B4, P_A25_B3, AND_A24_B4, Cout_A24_B3);

    wire AND_A25_B4;
    and and_a25_b4(AND_A25_B4, A[25], B[4]);
    wire P_A25_B4, Cout_A25_B4;
    full_adder add_a25_b4(P_A25_B4, Cout_A25_B4, P_A26_B3, AND_A25_B4, Cout_A25_B3);

    wire AND_A26_B4;
    and and_a26_b4(AND_A26_B4, A[26], B[4]);
    wire P_A26_B4, Cout_A26_B4;
    full_adder add_a26_b4(P_A26_B4, Cout_A26_B4, P_A27_B3, AND_A26_B4, Cout_A26_B3);

    wire AND_A27_B4;
    and and_a27_b4(AND_A27_B4, A[27], B[4]);
    wire P_A27_B4, Cout_A27_B4;
    full_adder add_a27_b4(P_A27_B4, Cout_A27_B4, P_A28_B3, AND_A27_B4, Cout_A27_B3);

    wire AND_A28_B4;
    and and_a28_b4(AND_A28_B4, A[28], B[4]);
    wire P_A28_B4, Cout_A28_B4;
    full_adder add_a28_b4(P_A28_B4, Cout_A28_B4, P_A29_B3, AND_A28_B4, Cout_A28_B3);

    wire AND_A29_B4;
    and and_a29_b4(AND_A29_B4, A[29], B[4]);
    wire P_A29_B4, Cout_A29_B4;
    full_adder add_a29_b4(P_A29_B4, Cout_A29_B4, P_A30_B3, AND_A29_B4, Cout_A29_B3);

    wire AND_A30_B4;
    and and_a30_b4(AND_A30_B4, A[30], B[4]);
    wire P_A30_B4, Cout_A30_B4;
    full_adder add_a30_b4(P_A30_B4, Cout_A30_B4, P_A31_B3, AND_A30_B4, Cout_A30_B3);

    wire AND_A31_B4;
    nand and_a31_b4(AND_A31_B4, A[31], B[4]);
    wire P_A31_B4, Cout_A31_B4;
    half_adder add_a31_b4(P_A31_B4, Cout_A31_B4, AND_A31_B4, Cout_A31_B3);

    wire AND_A0_B5;
    and and_a0_b5(AND_A0_B5, A[0], B[5]);
    wire P_A0_B5, Cout_A0_B5;
    full_adder add_a0_b5(P_A0_B5, Cout_A0_B5, P_A1_B4, AND_A0_B5, Cout_A0_B4);

    wire AND_A1_B5;
    and and_a1_b5(AND_A1_B5, A[1], B[5]);
    wire P_A1_B5, Cout_A1_B5;
    full_adder add_a1_b5(P_A1_B5, Cout_A1_B5, P_A2_B4, AND_A1_B5, Cout_A1_B4);

    wire AND_A2_B5;
    and and_a2_b5(AND_A2_B5, A[2], B[5]);
    wire P_A2_B5, Cout_A2_B5;
    full_adder add_a2_b5(P_A2_B5, Cout_A2_B5, P_A3_B4, AND_A2_B5, Cout_A2_B4);

    wire AND_A3_B5;
    and and_a3_b5(AND_A3_B5, A[3], B[5]);
    wire P_A3_B5, Cout_A3_B5;
    full_adder add_a3_b5(P_A3_B5, Cout_A3_B5, P_A4_B4, AND_A3_B5, Cout_A3_B4);

    wire AND_A4_B5;
    and and_a4_b5(AND_A4_B5, A[4], B[5]);
    wire P_A4_B5, Cout_A4_B5;
    full_adder add_a4_b5(P_A4_B5, Cout_A4_B5, P_A5_B4, AND_A4_B5, Cout_A4_B4);

    wire AND_A5_B5;
    and and_a5_b5(AND_A5_B5, A[5], B[5]);
    wire P_A5_B5, Cout_A5_B5;
    full_adder add_a5_b5(P_A5_B5, Cout_A5_B5, P_A6_B4, AND_A5_B5, Cout_A5_B4);

    wire AND_A6_B5;
    and and_a6_b5(AND_A6_B5, A[6], B[5]);
    wire P_A6_B5, Cout_A6_B5;
    full_adder add_a6_b5(P_A6_B5, Cout_A6_B5, P_A7_B4, AND_A6_B5, Cout_A6_B4);

    wire AND_A7_B5;
    and and_a7_b5(AND_A7_B5, A[7], B[5]);
    wire P_A7_B5, Cout_A7_B5;
    full_adder add_a7_b5(P_A7_B5, Cout_A7_B5, P_A8_B4, AND_A7_B5, Cout_A7_B4);

    wire AND_A8_B5;
    and and_a8_b5(AND_A8_B5, A[8], B[5]);
    wire P_A8_B5, Cout_A8_B5;
    full_adder add_a8_b5(P_A8_B5, Cout_A8_B5, P_A9_B4, AND_A8_B5, Cout_A8_B4);

    wire AND_A9_B5;
    and and_a9_b5(AND_A9_B5, A[9], B[5]);
    wire P_A9_B5, Cout_A9_B5;
    full_adder add_a9_b5(P_A9_B5, Cout_A9_B5, P_A10_B4, AND_A9_B5, Cout_A9_B4);

    wire AND_A10_B5;
    and and_a10_b5(AND_A10_B5, A[10], B[5]);
    wire P_A10_B5, Cout_A10_B5;
    full_adder add_a10_b5(P_A10_B5, Cout_A10_B5, P_A11_B4, AND_A10_B5, Cout_A10_B4);

    wire AND_A11_B5;
    and and_a11_b5(AND_A11_B5, A[11], B[5]);
    wire P_A11_B5, Cout_A11_B5;
    full_adder add_a11_b5(P_A11_B5, Cout_A11_B5, P_A12_B4, AND_A11_B5, Cout_A11_B4);

    wire AND_A12_B5;
    and and_a12_b5(AND_A12_B5, A[12], B[5]);
    wire P_A12_B5, Cout_A12_B5;
    full_adder add_a12_b5(P_A12_B5, Cout_A12_B5, P_A13_B4, AND_A12_B5, Cout_A12_B4);

    wire AND_A13_B5;
    and and_a13_b5(AND_A13_B5, A[13], B[5]);
    wire P_A13_B5, Cout_A13_B5;
    full_adder add_a13_b5(P_A13_B5, Cout_A13_B5, P_A14_B4, AND_A13_B5, Cout_A13_B4);

    wire AND_A14_B5;
    and and_a14_b5(AND_A14_B5, A[14], B[5]);
    wire P_A14_B5, Cout_A14_B5;
    full_adder add_a14_b5(P_A14_B5, Cout_A14_B5, P_A15_B4, AND_A14_B5, Cout_A14_B4);

    wire AND_A15_B5;
    and and_a15_b5(AND_A15_B5, A[15], B[5]);
    wire P_A15_B5, Cout_A15_B5;
    full_adder add_a15_b5(P_A15_B5, Cout_A15_B5, P_A16_B4, AND_A15_B5, Cout_A15_B4);

    wire AND_A16_B5;
    and and_a16_b5(AND_A16_B5, A[16], B[5]);
    wire P_A16_B5, Cout_A16_B5;
    full_adder add_a16_b5(P_A16_B5, Cout_A16_B5, P_A17_B4, AND_A16_B5, Cout_A16_B4);

    wire AND_A17_B5;
    and and_a17_b5(AND_A17_B5, A[17], B[5]);
    wire P_A17_B5, Cout_A17_B5;
    full_adder add_a17_b5(P_A17_B5, Cout_A17_B5, P_A18_B4, AND_A17_B5, Cout_A17_B4);

    wire AND_A18_B5;
    and and_a18_b5(AND_A18_B5, A[18], B[5]);
    wire P_A18_B5, Cout_A18_B5;
    full_adder add_a18_b5(P_A18_B5, Cout_A18_B5, P_A19_B4, AND_A18_B5, Cout_A18_B4);

    wire AND_A19_B5;
    and and_a19_b5(AND_A19_B5, A[19], B[5]);
    wire P_A19_B5, Cout_A19_B5;
    full_adder add_a19_b5(P_A19_B5, Cout_A19_B5, P_A20_B4, AND_A19_B5, Cout_A19_B4);

    wire AND_A20_B5;
    and and_a20_b5(AND_A20_B5, A[20], B[5]);
    wire P_A20_B5, Cout_A20_B5;
    full_adder add_a20_b5(P_A20_B5, Cout_A20_B5, P_A21_B4, AND_A20_B5, Cout_A20_B4);

    wire AND_A21_B5;
    and and_a21_b5(AND_A21_B5, A[21], B[5]);
    wire P_A21_B5, Cout_A21_B5;
    full_adder add_a21_b5(P_A21_B5, Cout_A21_B5, P_A22_B4, AND_A21_B5, Cout_A21_B4);

    wire AND_A22_B5;
    and and_a22_b5(AND_A22_B5, A[22], B[5]);
    wire P_A22_B5, Cout_A22_B5;
    full_adder add_a22_b5(P_A22_B5, Cout_A22_B5, P_A23_B4, AND_A22_B5, Cout_A22_B4);

    wire AND_A23_B5;
    and and_a23_b5(AND_A23_B5, A[23], B[5]);
    wire P_A23_B5, Cout_A23_B5;
    full_adder add_a23_b5(P_A23_B5, Cout_A23_B5, P_A24_B4, AND_A23_B5, Cout_A23_B4);

    wire AND_A24_B5;
    and and_a24_b5(AND_A24_B5, A[24], B[5]);
    wire P_A24_B5, Cout_A24_B5;
    full_adder add_a24_b5(P_A24_B5, Cout_A24_B5, P_A25_B4, AND_A24_B5, Cout_A24_B4);

    wire AND_A25_B5;
    and and_a25_b5(AND_A25_B5, A[25], B[5]);
    wire P_A25_B5, Cout_A25_B5;
    full_adder add_a25_b5(P_A25_B5, Cout_A25_B5, P_A26_B4, AND_A25_B5, Cout_A25_B4);

    wire AND_A26_B5;
    and and_a26_b5(AND_A26_B5, A[26], B[5]);
    wire P_A26_B5, Cout_A26_B5;
    full_adder add_a26_b5(P_A26_B5, Cout_A26_B5, P_A27_B4, AND_A26_B5, Cout_A26_B4);

    wire AND_A27_B5;
    and and_a27_b5(AND_A27_B5, A[27], B[5]);
    wire P_A27_B5, Cout_A27_B5;
    full_adder add_a27_b5(P_A27_B5, Cout_A27_B5, P_A28_B4, AND_A27_B5, Cout_A27_B4);

    wire AND_A28_B5;
    and and_a28_b5(AND_A28_B5, A[28], B[5]);
    wire P_A28_B5, Cout_A28_B5;
    full_adder add_a28_b5(P_A28_B5, Cout_A28_B5, P_A29_B4, AND_A28_B5, Cout_A28_B4);

    wire AND_A29_B5;
    and and_a29_b5(AND_A29_B5, A[29], B[5]);
    wire P_A29_B5, Cout_A29_B5;
    full_adder add_a29_b5(P_A29_B5, Cout_A29_B5, P_A30_B4, AND_A29_B5, Cout_A29_B4);

    wire AND_A30_B5;
    and and_a30_b5(AND_A30_B5, A[30], B[5]);
    wire P_A30_B5, Cout_A30_B5;
    full_adder add_a30_b5(P_A30_B5, Cout_A30_B5, P_A31_B4, AND_A30_B5, Cout_A30_B4);

    wire AND_A31_B5;
    nand and_a31_b5(AND_A31_B5, A[31], B[5]);
    wire P_A31_B5, Cout_A31_B5;
    half_adder add_a31_b5(P_A31_B5, Cout_A31_B5, AND_A31_B5, Cout_A31_B4);

    wire AND_A0_B6;
    and and_a0_b6(AND_A0_B6, A[0], B[6]);
    wire P_A0_B6, Cout_A0_B6;
    full_adder add_a0_b6(P_A0_B6, Cout_A0_B6, P_A1_B5, AND_A0_B6, Cout_A0_B5);

    wire AND_A1_B6;
    and and_a1_b6(AND_A1_B6, A[1], B[6]);
    wire P_A1_B6, Cout_A1_B6;
    full_adder add_a1_b6(P_A1_B6, Cout_A1_B6, P_A2_B5, AND_A1_B6, Cout_A1_B5);

    wire AND_A2_B6;
    and and_a2_b6(AND_A2_B6, A[2], B[6]);
    wire P_A2_B6, Cout_A2_B6;
    full_adder add_a2_b6(P_A2_B6, Cout_A2_B6, P_A3_B5, AND_A2_B6, Cout_A2_B5);

    wire AND_A3_B6;
    and and_a3_b6(AND_A3_B6, A[3], B[6]);
    wire P_A3_B6, Cout_A3_B6;
    full_adder add_a3_b6(P_A3_B6, Cout_A3_B6, P_A4_B5, AND_A3_B6, Cout_A3_B5);

    wire AND_A4_B6;
    and and_a4_b6(AND_A4_B6, A[4], B[6]);
    wire P_A4_B6, Cout_A4_B6;
    full_adder add_a4_b6(P_A4_B6, Cout_A4_B6, P_A5_B5, AND_A4_B6, Cout_A4_B5);

    wire AND_A5_B6;
    and and_a5_b6(AND_A5_B6, A[5], B[6]);
    wire P_A5_B6, Cout_A5_B6;
    full_adder add_a5_b6(P_A5_B6, Cout_A5_B6, P_A6_B5, AND_A5_B6, Cout_A5_B5);

    wire AND_A6_B6;
    and and_a6_b6(AND_A6_B6, A[6], B[6]);
    wire P_A6_B6, Cout_A6_B6;
    full_adder add_a6_b6(P_A6_B6, Cout_A6_B6, P_A7_B5, AND_A6_B6, Cout_A6_B5);

    wire AND_A7_B6;
    and and_a7_b6(AND_A7_B6, A[7], B[6]);
    wire P_A7_B6, Cout_A7_B6;
    full_adder add_a7_b6(P_A7_B6, Cout_A7_B6, P_A8_B5, AND_A7_B6, Cout_A7_B5);

    wire AND_A8_B6;
    and and_a8_b6(AND_A8_B6, A[8], B[6]);
    wire P_A8_B6, Cout_A8_B6;
    full_adder add_a8_b6(P_A8_B6, Cout_A8_B6, P_A9_B5, AND_A8_B6, Cout_A8_B5);

    wire AND_A9_B6;
    and and_a9_b6(AND_A9_B6, A[9], B[6]);
    wire P_A9_B6, Cout_A9_B6;
    full_adder add_a9_b6(P_A9_B6, Cout_A9_B6, P_A10_B5, AND_A9_B6, Cout_A9_B5);

    wire AND_A10_B6;
    and and_a10_b6(AND_A10_B6, A[10], B[6]);
    wire P_A10_B6, Cout_A10_B6;
    full_adder add_a10_b6(P_A10_B6, Cout_A10_B6, P_A11_B5, AND_A10_B6, Cout_A10_B5);

    wire AND_A11_B6;
    and and_a11_b6(AND_A11_B6, A[11], B[6]);
    wire P_A11_B6, Cout_A11_B6;
    full_adder add_a11_b6(P_A11_B6, Cout_A11_B6, P_A12_B5, AND_A11_B6, Cout_A11_B5);

    wire AND_A12_B6;
    and and_a12_b6(AND_A12_B6, A[12], B[6]);
    wire P_A12_B6, Cout_A12_B6;
    full_adder add_a12_b6(P_A12_B6, Cout_A12_B6, P_A13_B5, AND_A12_B6, Cout_A12_B5);

    wire AND_A13_B6;
    and and_a13_b6(AND_A13_B6, A[13], B[6]);
    wire P_A13_B6, Cout_A13_B6;
    full_adder add_a13_b6(P_A13_B6, Cout_A13_B6, P_A14_B5, AND_A13_B6, Cout_A13_B5);

    wire AND_A14_B6;
    and and_a14_b6(AND_A14_B6, A[14], B[6]);
    wire P_A14_B6, Cout_A14_B6;
    full_adder add_a14_b6(P_A14_B6, Cout_A14_B6, P_A15_B5, AND_A14_B6, Cout_A14_B5);

    wire AND_A15_B6;
    and and_a15_b6(AND_A15_B6, A[15], B[6]);
    wire P_A15_B6, Cout_A15_B6;
    full_adder add_a15_b6(P_A15_B6, Cout_A15_B6, P_A16_B5, AND_A15_B6, Cout_A15_B5);

    wire AND_A16_B6;
    and and_a16_b6(AND_A16_B6, A[16], B[6]);
    wire P_A16_B6, Cout_A16_B6;
    full_adder add_a16_b6(P_A16_B6, Cout_A16_B6, P_A17_B5, AND_A16_B6, Cout_A16_B5);

    wire AND_A17_B6;
    and and_a17_b6(AND_A17_B6, A[17], B[6]);
    wire P_A17_B6, Cout_A17_B6;
    full_adder add_a17_b6(P_A17_B6, Cout_A17_B6, P_A18_B5, AND_A17_B6, Cout_A17_B5);

    wire AND_A18_B6;
    and and_a18_b6(AND_A18_B6, A[18], B[6]);
    wire P_A18_B6, Cout_A18_B6;
    full_adder add_a18_b6(P_A18_B6, Cout_A18_B6, P_A19_B5, AND_A18_B6, Cout_A18_B5);

    wire AND_A19_B6;
    and and_a19_b6(AND_A19_B6, A[19], B[6]);
    wire P_A19_B6, Cout_A19_B6;
    full_adder add_a19_b6(P_A19_B6, Cout_A19_B6, P_A20_B5, AND_A19_B6, Cout_A19_B5);

    wire AND_A20_B6;
    and and_a20_b6(AND_A20_B6, A[20], B[6]);
    wire P_A20_B6, Cout_A20_B6;
    full_adder add_a20_b6(P_A20_B6, Cout_A20_B6, P_A21_B5, AND_A20_B6, Cout_A20_B5);

    wire AND_A21_B6;
    and and_a21_b6(AND_A21_B6, A[21], B[6]);
    wire P_A21_B6, Cout_A21_B6;
    full_adder add_a21_b6(P_A21_B6, Cout_A21_B6, P_A22_B5, AND_A21_B6, Cout_A21_B5);

    wire AND_A22_B6;
    and and_a22_b6(AND_A22_B6, A[22], B[6]);
    wire P_A22_B6, Cout_A22_B6;
    full_adder add_a22_b6(P_A22_B6, Cout_A22_B6, P_A23_B5, AND_A22_B6, Cout_A22_B5);

    wire AND_A23_B6;
    and and_a23_b6(AND_A23_B6, A[23], B[6]);
    wire P_A23_B6, Cout_A23_B6;
    full_adder add_a23_b6(P_A23_B6, Cout_A23_B6, P_A24_B5, AND_A23_B6, Cout_A23_B5);

    wire AND_A24_B6;
    and and_a24_b6(AND_A24_B6, A[24], B[6]);
    wire P_A24_B6, Cout_A24_B6;
    full_adder add_a24_b6(P_A24_B6, Cout_A24_B6, P_A25_B5, AND_A24_B6, Cout_A24_B5);

    wire AND_A25_B6;
    and and_a25_b6(AND_A25_B6, A[25], B[6]);
    wire P_A25_B6, Cout_A25_B6;
    full_adder add_a25_b6(P_A25_B6, Cout_A25_B6, P_A26_B5, AND_A25_B6, Cout_A25_B5);

    wire AND_A26_B6;
    and and_a26_b6(AND_A26_B6, A[26], B[6]);
    wire P_A26_B6, Cout_A26_B6;
    full_adder add_a26_b6(P_A26_B6, Cout_A26_B6, P_A27_B5, AND_A26_B6, Cout_A26_B5);

    wire AND_A27_B6;
    and and_a27_b6(AND_A27_B6, A[27], B[6]);
    wire P_A27_B6, Cout_A27_B6;
    full_adder add_a27_b6(P_A27_B6, Cout_A27_B6, P_A28_B5, AND_A27_B6, Cout_A27_B5);

    wire AND_A28_B6;
    and and_a28_b6(AND_A28_B6, A[28], B[6]);
    wire P_A28_B6, Cout_A28_B6;
    full_adder add_a28_b6(P_A28_B6, Cout_A28_B6, P_A29_B5, AND_A28_B6, Cout_A28_B5);

    wire AND_A29_B6;
    and and_a29_b6(AND_A29_B6, A[29], B[6]);
    wire P_A29_B6, Cout_A29_B6;
    full_adder add_a29_b6(P_A29_B6, Cout_A29_B6, P_A30_B5, AND_A29_B6, Cout_A29_B5);

    wire AND_A30_B6;
    and and_a30_b6(AND_A30_B6, A[30], B[6]);
    wire P_A30_B6, Cout_A30_B6;
    full_adder add_a30_b6(P_A30_B6, Cout_A30_B6, P_A31_B5, AND_A30_B6, Cout_A30_B5);

    wire AND_A31_B6;
    nand and_a31_b6(AND_A31_B6, A[31], B[6]);
    wire P_A31_B6, Cout_A31_B6;
    half_adder add_a31_b6(P_A31_B6, Cout_A31_B6, AND_A31_B6, Cout_A31_B5);

    wire AND_A0_B7;
    and and_a0_b7(AND_A0_B7, A[0], B[7]);
    wire P_A0_B7, Cout_A0_B7;
    full_adder add_a0_b7(P_A0_B7, Cout_A0_B7, P_A1_B6, AND_A0_B7, Cout_A0_B6);

    wire AND_A1_B7;
    and and_a1_b7(AND_A1_B7, A[1], B[7]);
    wire P_A1_B7, Cout_A1_B7;
    full_adder add_a1_b7(P_A1_B7, Cout_A1_B7, P_A2_B6, AND_A1_B7, Cout_A1_B6);

    wire AND_A2_B7;
    and and_a2_b7(AND_A2_B7, A[2], B[7]);
    wire P_A2_B7, Cout_A2_B7;
    full_adder add_a2_b7(P_A2_B7, Cout_A2_B7, P_A3_B6, AND_A2_B7, Cout_A2_B6);

    wire AND_A3_B7;
    and and_a3_b7(AND_A3_B7, A[3], B[7]);
    wire P_A3_B7, Cout_A3_B7;
    full_adder add_a3_b7(P_A3_B7, Cout_A3_B7, P_A4_B6, AND_A3_B7, Cout_A3_B6);

    wire AND_A4_B7;
    and and_a4_b7(AND_A4_B7, A[4], B[7]);
    wire P_A4_B7, Cout_A4_B7;
    full_adder add_a4_b7(P_A4_B7, Cout_A4_B7, P_A5_B6, AND_A4_B7, Cout_A4_B6);

    wire AND_A5_B7;
    and and_a5_b7(AND_A5_B7, A[5], B[7]);
    wire P_A5_B7, Cout_A5_B7;
    full_adder add_a5_b7(P_A5_B7, Cout_A5_B7, P_A6_B6, AND_A5_B7, Cout_A5_B6);

    wire AND_A6_B7;
    and and_a6_b7(AND_A6_B7, A[6], B[7]);
    wire P_A6_B7, Cout_A6_B7;
    full_adder add_a6_b7(P_A6_B7, Cout_A6_B7, P_A7_B6, AND_A6_B7, Cout_A6_B6);

    wire AND_A7_B7;
    and and_a7_b7(AND_A7_B7, A[7], B[7]);
    wire P_A7_B7, Cout_A7_B7;
    full_adder add_a7_b7(P_A7_B7, Cout_A7_B7, P_A8_B6, AND_A7_B7, Cout_A7_B6);

    wire AND_A8_B7;
    and and_a8_b7(AND_A8_B7, A[8], B[7]);
    wire P_A8_B7, Cout_A8_B7;
    full_adder add_a8_b7(P_A8_B7, Cout_A8_B7, P_A9_B6, AND_A8_B7, Cout_A8_B6);

    wire AND_A9_B7;
    and and_a9_b7(AND_A9_B7, A[9], B[7]);
    wire P_A9_B7, Cout_A9_B7;
    full_adder add_a9_b7(P_A9_B7, Cout_A9_B7, P_A10_B6, AND_A9_B7, Cout_A9_B6);

    wire AND_A10_B7;
    and and_a10_b7(AND_A10_B7, A[10], B[7]);
    wire P_A10_B7, Cout_A10_B7;
    full_adder add_a10_b7(P_A10_B7, Cout_A10_B7, P_A11_B6, AND_A10_B7, Cout_A10_B6);

    wire AND_A11_B7;
    and and_a11_b7(AND_A11_B7, A[11], B[7]);
    wire P_A11_B7, Cout_A11_B7;
    full_adder add_a11_b7(P_A11_B7, Cout_A11_B7, P_A12_B6, AND_A11_B7, Cout_A11_B6);

    wire AND_A12_B7;
    and and_a12_b7(AND_A12_B7, A[12], B[7]);
    wire P_A12_B7, Cout_A12_B7;
    full_adder add_a12_b7(P_A12_B7, Cout_A12_B7, P_A13_B6, AND_A12_B7, Cout_A12_B6);

    wire AND_A13_B7;
    and and_a13_b7(AND_A13_B7, A[13], B[7]);
    wire P_A13_B7, Cout_A13_B7;
    full_adder add_a13_b7(P_A13_B7, Cout_A13_B7, P_A14_B6, AND_A13_B7, Cout_A13_B6);

    wire AND_A14_B7;
    and and_a14_b7(AND_A14_B7, A[14], B[7]);
    wire P_A14_B7, Cout_A14_B7;
    full_adder add_a14_b7(P_A14_B7, Cout_A14_B7, P_A15_B6, AND_A14_B7, Cout_A14_B6);

    wire AND_A15_B7;
    and and_a15_b7(AND_A15_B7, A[15], B[7]);
    wire P_A15_B7, Cout_A15_B7;
    full_adder add_a15_b7(P_A15_B7, Cout_A15_B7, P_A16_B6, AND_A15_B7, Cout_A15_B6);

    wire AND_A16_B7;
    and and_a16_b7(AND_A16_B7, A[16], B[7]);
    wire P_A16_B7, Cout_A16_B7;
    full_adder add_a16_b7(P_A16_B7, Cout_A16_B7, P_A17_B6, AND_A16_B7, Cout_A16_B6);

    wire AND_A17_B7;
    and and_a17_b7(AND_A17_B7, A[17], B[7]);
    wire P_A17_B7, Cout_A17_B7;
    full_adder add_a17_b7(P_A17_B7, Cout_A17_B7, P_A18_B6, AND_A17_B7, Cout_A17_B6);

    wire AND_A18_B7;
    and and_a18_b7(AND_A18_B7, A[18], B[7]);
    wire P_A18_B7, Cout_A18_B7;
    full_adder add_a18_b7(P_A18_B7, Cout_A18_B7, P_A19_B6, AND_A18_B7, Cout_A18_B6);

    wire AND_A19_B7;
    and and_a19_b7(AND_A19_B7, A[19], B[7]);
    wire P_A19_B7, Cout_A19_B7;
    full_adder add_a19_b7(P_A19_B7, Cout_A19_B7, P_A20_B6, AND_A19_B7, Cout_A19_B6);

    wire AND_A20_B7;
    and and_a20_b7(AND_A20_B7, A[20], B[7]);
    wire P_A20_B7, Cout_A20_B7;
    full_adder add_a20_b7(P_A20_B7, Cout_A20_B7, P_A21_B6, AND_A20_B7, Cout_A20_B6);

    wire AND_A21_B7;
    and and_a21_b7(AND_A21_B7, A[21], B[7]);
    wire P_A21_B7, Cout_A21_B7;
    full_adder add_a21_b7(P_A21_B7, Cout_A21_B7, P_A22_B6, AND_A21_B7, Cout_A21_B6);

    wire AND_A22_B7;
    and and_a22_b7(AND_A22_B7, A[22], B[7]);
    wire P_A22_B7, Cout_A22_B7;
    full_adder add_a22_b7(P_A22_B7, Cout_A22_B7, P_A23_B6, AND_A22_B7, Cout_A22_B6);

    wire AND_A23_B7;
    and and_a23_b7(AND_A23_B7, A[23], B[7]);
    wire P_A23_B7, Cout_A23_B7;
    full_adder add_a23_b7(P_A23_B7, Cout_A23_B7, P_A24_B6, AND_A23_B7, Cout_A23_B6);

    wire AND_A24_B7;
    and and_a24_b7(AND_A24_B7, A[24], B[7]);
    wire P_A24_B7, Cout_A24_B7;
    full_adder add_a24_b7(P_A24_B7, Cout_A24_B7, P_A25_B6, AND_A24_B7, Cout_A24_B6);

    wire AND_A25_B7;
    and and_a25_b7(AND_A25_B7, A[25], B[7]);
    wire P_A25_B7, Cout_A25_B7;
    full_adder add_a25_b7(P_A25_B7, Cout_A25_B7, P_A26_B6, AND_A25_B7, Cout_A25_B6);

    wire AND_A26_B7;
    and and_a26_b7(AND_A26_B7, A[26], B[7]);
    wire P_A26_B7, Cout_A26_B7;
    full_adder add_a26_b7(P_A26_B7, Cout_A26_B7, P_A27_B6, AND_A26_B7, Cout_A26_B6);

    wire AND_A27_B7;
    and and_a27_b7(AND_A27_B7, A[27], B[7]);
    wire P_A27_B7, Cout_A27_B7;
    full_adder add_a27_b7(P_A27_B7, Cout_A27_B7, P_A28_B6, AND_A27_B7, Cout_A27_B6);

    wire AND_A28_B7;
    and and_a28_b7(AND_A28_B7, A[28], B[7]);
    wire P_A28_B7, Cout_A28_B7;
    full_adder add_a28_b7(P_A28_B7, Cout_A28_B7, P_A29_B6, AND_A28_B7, Cout_A28_B6);

    wire AND_A29_B7;
    and and_a29_b7(AND_A29_B7, A[29], B[7]);
    wire P_A29_B7, Cout_A29_B7;
    full_adder add_a29_b7(P_A29_B7, Cout_A29_B7, P_A30_B6, AND_A29_B7, Cout_A29_B6);

    wire AND_A30_B7;
    and and_a30_b7(AND_A30_B7, A[30], B[7]);
    wire P_A30_B7, Cout_A30_B7;
    full_adder add_a30_b7(P_A30_B7, Cout_A30_B7, P_A31_B6, AND_A30_B7, Cout_A30_B6);

    wire AND_A31_B7;
    nand and_a31_b7(AND_A31_B7, A[31], B[7]);
    wire P_A31_B7, Cout_A31_B7;
    half_adder add_a31_b7(P_A31_B7, Cout_A31_B7, AND_A31_B7, Cout_A31_B6);

    wire AND_A0_B8;
    and and_a0_b8(AND_A0_B8, A[0], B[8]);
    wire P_A0_B8, Cout_A0_B8;
    full_adder add_a0_b8(P_A0_B8, Cout_A0_B8, P_A1_B7, AND_A0_B8, Cout_A0_B7);

    wire AND_A1_B8;
    and and_a1_b8(AND_A1_B8, A[1], B[8]);
    wire P_A1_B8, Cout_A1_B8;
    full_adder add_a1_b8(P_A1_B8, Cout_A1_B8, P_A2_B7, AND_A1_B8, Cout_A1_B7);

    wire AND_A2_B8;
    and and_a2_b8(AND_A2_B8, A[2], B[8]);
    wire P_A2_B8, Cout_A2_B8;
    full_adder add_a2_b8(P_A2_B8, Cout_A2_B8, P_A3_B7, AND_A2_B8, Cout_A2_B7);

    wire AND_A3_B8;
    and and_a3_b8(AND_A3_B8, A[3], B[8]);
    wire P_A3_B8, Cout_A3_B8;
    full_adder add_a3_b8(P_A3_B8, Cout_A3_B8, P_A4_B7, AND_A3_B8, Cout_A3_B7);

    wire AND_A4_B8;
    and and_a4_b8(AND_A4_B8, A[4], B[8]);
    wire P_A4_B8, Cout_A4_B8;
    full_adder add_a4_b8(P_A4_B8, Cout_A4_B8, P_A5_B7, AND_A4_B8, Cout_A4_B7);

    wire AND_A5_B8;
    and and_a5_b8(AND_A5_B8, A[5], B[8]);
    wire P_A5_B8, Cout_A5_B8;
    full_adder add_a5_b8(P_A5_B8, Cout_A5_B8, P_A6_B7, AND_A5_B8, Cout_A5_B7);

    wire AND_A6_B8;
    and and_a6_b8(AND_A6_B8, A[6], B[8]);
    wire P_A6_B8, Cout_A6_B8;
    full_adder add_a6_b8(P_A6_B8, Cout_A6_B8, P_A7_B7, AND_A6_B8, Cout_A6_B7);

    wire AND_A7_B8;
    and and_a7_b8(AND_A7_B8, A[7], B[8]);
    wire P_A7_B8, Cout_A7_B8;
    full_adder add_a7_b8(P_A7_B8, Cout_A7_B8, P_A8_B7, AND_A7_B8, Cout_A7_B7);

    wire AND_A8_B8;
    and and_a8_b8(AND_A8_B8, A[8], B[8]);
    wire P_A8_B8, Cout_A8_B8;
    full_adder add_a8_b8(P_A8_B8, Cout_A8_B8, P_A9_B7, AND_A8_B8, Cout_A8_B7);

    wire AND_A9_B8;
    and and_a9_b8(AND_A9_B8, A[9], B[8]);
    wire P_A9_B8, Cout_A9_B8;
    full_adder add_a9_b8(P_A9_B8, Cout_A9_B8, P_A10_B7, AND_A9_B8, Cout_A9_B7);

    wire AND_A10_B8;
    and and_a10_b8(AND_A10_B8, A[10], B[8]);
    wire P_A10_B8, Cout_A10_B8;
    full_adder add_a10_b8(P_A10_B8, Cout_A10_B8, P_A11_B7, AND_A10_B8, Cout_A10_B7);

    wire AND_A11_B8;
    and and_a11_b8(AND_A11_B8, A[11], B[8]);
    wire P_A11_B8, Cout_A11_B8;
    full_adder add_a11_b8(P_A11_B8, Cout_A11_B8, P_A12_B7, AND_A11_B8, Cout_A11_B7);

    wire AND_A12_B8;
    and and_a12_b8(AND_A12_B8, A[12], B[8]);
    wire P_A12_B8, Cout_A12_B8;
    full_adder add_a12_b8(P_A12_B8, Cout_A12_B8, P_A13_B7, AND_A12_B8, Cout_A12_B7);

    wire AND_A13_B8;
    and and_a13_b8(AND_A13_B8, A[13], B[8]);
    wire P_A13_B8, Cout_A13_B8;
    full_adder add_a13_b8(P_A13_B8, Cout_A13_B8, P_A14_B7, AND_A13_B8, Cout_A13_B7);

    wire AND_A14_B8;
    and and_a14_b8(AND_A14_B8, A[14], B[8]);
    wire P_A14_B8, Cout_A14_B8;
    full_adder add_a14_b8(P_A14_B8, Cout_A14_B8, P_A15_B7, AND_A14_B8, Cout_A14_B7);

    wire AND_A15_B8;
    and and_a15_b8(AND_A15_B8, A[15], B[8]);
    wire P_A15_B8, Cout_A15_B8;
    full_adder add_a15_b8(P_A15_B8, Cout_A15_B8, P_A16_B7, AND_A15_B8, Cout_A15_B7);

    wire AND_A16_B8;
    and and_a16_b8(AND_A16_B8, A[16], B[8]);
    wire P_A16_B8, Cout_A16_B8;
    full_adder add_a16_b8(P_A16_B8, Cout_A16_B8, P_A17_B7, AND_A16_B8, Cout_A16_B7);

    wire AND_A17_B8;
    and and_a17_b8(AND_A17_B8, A[17], B[8]);
    wire P_A17_B8, Cout_A17_B8;
    full_adder add_a17_b8(P_A17_B8, Cout_A17_B8, P_A18_B7, AND_A17_B8, Cout_A17_B7);

    wire AND_A18_B8;
    and and_a18_b8(AND_A18_B8, A[18], B[8]);
    wire P_A18_B8, Cout_A18_B8;
    full_adder add_a18_b8(P_A18_B8, Cout_A18_B8, P_A19_B7, AND_A18_B8, Cout_A18_B7);

    wire AND_A19_B8;
    and and_a19_b8(AND_A19_B8, A[19], B[8]);
    wire P_A19_B8, Cout_A19_B8;
    full_adder add_a19_b8(P_A19_B8, Cout_A19_B8, P_A20_B7, AND_A19_B8, Cout_A19_B7);

    wire AND_A20_B8;
    and and_a20_b8(AND_A20_B8, A[20], B[8]);
    wire P_A20_B8, Cout_A20_B8;
    full_adder add_a20_b8(P_A20_B8, Cout_A20_B8, P_A21_B7, AND_A20_B8, Cout_A20_B7);

    wire AND_A21_B8;
    and and_a21_b8(AND_A21_B8, A[21], B[8]);
    wire P_A21_B8, Cout_A21_B8;
    full_adder add_a21_b8(P_A21_B8, Cout_A21_B8, P_A22_B7, AND_A21_B8, Cout_A21_B7);

    wire AND_A22_B8;
    and and_a22_b8(AND_A22_B8, A[22], B[8]);
    wire P_A22_B8, Cout_A22_B8;
    full_adder add_a22_b8(P_A22_B8, Cout_A22_B8, P_A23_B7, AND_A22_B8, Cout_A22_B7);

    wire AND_A23_B8;
    and and_a23_b8(AND_A23_B8, A[23], B[8]);
    wire P_A23_B8, Cout_A23_B8;
    full_adder add_a23_b8(P_A23_B8, Cout_A23_B8, P_A24_B7, AND_A23_B8, Cout_A23_B7);

    wire AND_A24_B8;
    and and_a24_b8(AND_A24_B8, A[24], B[8]);
    wire P_A24_B8, Cout_A24_B8;
    full_adder add_a24_b8(P_A24_B8, Cout_A24_B8, P_A25_B7, AND_A24_B8, Cout_A24_B7);

    wire AND_A25_B8;
    and and_a25_b8(AND_A25_B8, A[25], B[8]);
    wire P_A25_B8, Cout_A25_B8;
    full_adder add_a25_b8(P_A25_B8, Cout_A25_B8, P_A26_B7, AND_A25_B8, Cout_A25_B7);

    wire AND_A26_B8;
    and and_a26_b8(AND_A26_B8, A[26], B[8]);
    wire P_A26_B8, Cout_A26_B8;
    full_adder add_a26_b8(P_A26_B8, Cout_A26_B8, P_A27_B7, AND_A26_B8, Cout_A26_B7);

    wire AND_A27_B8;
    and and_a27_b8(AND_A27_B8, A[27], B[8]);
    wire P_A27_B8, Cout_A27_B8;
    full_adder add_a27_b8(P_A27_B8, Cout_A27_B8, P_A28_B7, AND_A27_B8, Cout_A27_B7);

    wire AND_A28_B8;
    and and_a28_b8(AND_A28_B8, A[28], B[8]);
    wire P_A28_B8, Cout_A28_B8;
    full_adder add_a28_b8(P_A28_B8, Cout_A28_B8, P_A29_B7, AND_A28_B8, Cout_A28_B7);

    wire AND_A29_B8;
    and and_a29_b8(AND_A29_B8, A[29], B[8]);
    wire P_A29_B8, Cout_A29_B8;
    full_adder add_a29_b8(P_A29_B8, Cout_A29_B8, P_A30_B7, AND_A29_B8, Cout_A29_B7);

    wire AND_A30_B8;
    and and_a30_b8(AND_A30_B8, A[30], B[8]);
    wire P_A30_B8, Cout_A30_B8;
    full_adder add_a30_b8(P_A30_B8, Cout_A30_B8, P_A31_B7, AND_A30_B8, Cout_A30_B7);

    wire AND_A31_B8;
    nand and_a31_b8(AND_A31_B8, A[31], B[8]);
    wire P_A31_B8, Cout_A31_B8;
    half_adder add_a31_b8(P_A31_B8, Cout_A31_B8, AND_A31_B8, Cout_A31_B7);

    wire AND_A0_B9;
    and and_a0_b9(AND_A0_B9, A[0], B[9]);
    wire P_A0_B9, Cout_A0_B9;
    full_adder add_a0_b9(P_A0_B9, Cout_A0_B9, P_A1_B8, AND_A0_B9, Cout_A0_B8);

    wire AND_A1_B9;
    and and_a1_b9(AND_A1_B9, A[1], B[9]);
    wire P_A1_B9, Cout_A1_B9;
    full_adder add_a1_b9(P_A1_B9, Cout_A1_B9, P_A2_B8, AND_A1_B9, Cout_A1_B8);

    wire AND_A2_B9;
    and and_a2_b9(AND_A2_B9, A[2], B[9]);
    wire P_A2_B9, Cout_A2_B9;
    full_adder add_a2_b9(P_A2_B9, Cout_A2_B9, P_A3_B8, AND_A2_B9, Cout_A2_B8);

    wire AND_A3_B9;
    and and_a3_b9(AND_A3_B9, A[3], B[9]);
    wire P_A3_B9, Cout_A3_B9;
    full_adder add_a3_b9(P_A3_B9, Cout_A3_B9, P_A4_B8, AND_A3_B9, Cout_A3_B8);

    wire AND_A4_B9;
    and and_a4_b9(AND_A4_B9, A[4], B[9]);
    wire P_A4_B9, Cout_A4_B9;
    full_adder add_a4_b9(P_A4_B9, Cout_A4_B9, P_A5_B8, AND_A4_B9, Cout_A4_B8);

    wire AND_A5_B9;
    and and_a5_b9(AND_A5_B9, A[5], B[9]);
    wire P_A5_B9, Cout_A5_B9;
    full_adder add_a5_b9(P_A5_B9, Cout_A5_B9, P_A6_B8, AND_A5_B9, Cout_A5_B8);

    wire AND_A6_B9;
    and and_a6_b9(AND_A6_B9, A[6], B[9]);
    wire P_A6_B9, Cout_A6_B9;
    full_adder add_a6_b9(P_A6_B9, Cout_A6_B9, P_A7_B8, AND_A6_B9, Cout_A6_B8);

    wire AND_A7_B9;
    and and_a7_b9(AND_A7_B9, A[7], B[9]);
    wire P_A7_B9, Cout_A7_B9;
    full_adder add_a7_b9(P_A7_B9, Cout_A7_B9, P_A8_B8, AND_A7_B9, Cout_A7_B8);

    wire AND_A8_B9;
    and and_a8_b9(AND_A8_B9, A[8], B[9]);
    wire P_A8_B9, Cout_A8_B9;
    full_adder add_a8_b9(P_A8_B9, Cout_A8_B9, P_A9_B8, AND_A8_B9, Cout_A8_B8);

    wire AND_A9_B9;
    and and_a9_b9(AND_A9_B9, A[9], B[9]);
    wire P_A9_B9, Cout_A9_B9;
    full_adder add_a9_b9(P_A9_B9, Cout_A9_B9, P_A10_B8, AND_A9_B9, Cout_A9_B8);

    wire AND_A10_B9;
    and and_a10_b9(AND_A10_B9, A[10], B[9]);
    wire P_A10_B9, Cout_A10_B9;
    full_adder add_a10_b9(P_A10_B9, Cout_A10_B9, P_A11_B8, AND_A10_B9, Cout_A10_B8);

    wire AND_A11_B9;
    and and_a11_b9(AND_A11_B9, A[11], B[9]);
    wire P_A11_B9, Cout_A11_B9;
    full_adder add_a11_b9(P_A11_B9, Cout_A11_B9, P_A12_B8, AND_A11_B9, Cout_A11_B8);

    wire AND_A12_B9;
    and and_a12_b9(AND_A12_B9, A[12], B[9]);
    wire P_A12_B9, Cout_A12_B9;
    full_adder add_a12_b9(P_A12_B9, Cout_A12_B9, P_A13_B8, AND_A12_B9, Cout_A12_B8);

    wire AND_A13_B9;
    and and_a13_b9(AND_A13_B9, A[13], B[9]);
    wire P_A13_B9, Cout_A13_B9;
    full_adder add_a13_b9(P_A13_B9, Cout_A13_B9, P_A14_B8, AND_A13_B9, Cout_A13_B8);

    wire AND_A14_B9;
    and and_a14_b9(AND_A14_B9, A[14], B[9]);
    wire P_A14_B9, Cout_A14_B9;
    full_adder add_a14_b9(P_A14_B9, Cout_A14_B9, P_A15_B8, AND_A14_B9, Cout_A14_B8);

    wire AND_A15_B9;
    and and_a15_b9(AND_A15_B9, A[15], B[9]);
    wire P_A15_B9, Cout_A15_B9;
    full_adder add_a15_b9(P_A15_B9, Cout_A15_B9, P_A16_B8, AND_A15_B9, Cout_A15_B8);

    wire AND_A16_B9;
    and and_a16_b9(AND_A16_B9, A[16], B[9]);
    wire P_A16_B9, Cout_A16_B9;
    full_adder add_a16_b9(P_A16_B9, Cout_A16_B9, P_A17_B8, AND_A16_B9, Cout_A16_B8);

    wire AND_A17_B9;
    and and_a17_b9(AND_A17_B9, A[17], B[9]);
    wire P_A17_B9, Cout_A17_B9;
    full_adder add_a17_b9(P_A17_B9, Cout_A17_B9, P_A18_B8, AND_A17_B9, Cout_A17_B8);

    wire AND_A18_B9;
    and and_a18_b9(AND_A18_B9, A[18], B[9]);
    wire P_A18_B9, Cout_A18_B9;
    full_adder add_a18_b9(P_A18_B9, Cout_A18_B9, P_A19_B8, AND_A18_B9, Cout_A18_B8);

    wire AND_A19_B9;
    and and_a19_b9(AND_A19_B9, A[19], B[9]);
    wire P_A19_B9, Cout_A19_B9;
    full_adder add_a19_b9(P_A19_B9, Cout_A19_B9, P_A20_B8, AND_A19_B9, Cout_A19_B8);

    wire AND_A20_B9;
    and and_a20_b9(AND_A20_B9, A[20], B[9]);
    wire P_A20_B9, Cout_A20_B9;
    full_adder add_a20_b9(P_A20_B9, Cout_A20_B9, P_A21_B8, AND_A20_B9, Cout_A20_B8);

    wire AND_A21_B9;
    and and_a21_b9(AND_A21_B9, A[21], B[9]);
    wire P_A21_B9, Cout_A21_B9;
    full_adder add_a21_b9(P_A21_B9, Cout_A21_B9, P_A22_B8, AND_A21_B9, Cout_A21_B8);

    wire AND_A22_B9;
    and and_a22_b9(AND_A22_B9, A[22], B[9]);
    wire P_A22_B9, Cout_A22_B9;
    full_adder add_a22_b9(P_A22_B9, Cout_A22_B9, P_A23_B8, AND_A22_B9, Cout_A22_B8);

    wire AND_A23_B9;
    and and_a23_b9(AND_A23_B9, A[23], B[9]);
    wire P_A23_B9, Cout_A23_B9;
    full_adder add_a23_b9(P_A23_B9, Cout_A23_B9, P_A24_B8, AND_A23_B9, Cout_A23_B8);

    wire AND_A24_B9;
    and and_a24_b9(AND_A24_B9, A[24], B[9]);
    wire P_A24_B9, Cout_A24_B9;
    full_adder add_a24_b9(P_A24_B9, Cout_A24_B9, P_A25_B8, AND_A24_B9, Cout_A24_B8);

    wire AND_A25_B9;
    and and_a25_b9(AND_A25_B9, A[25], B[9]);
    wire P_A25_B9, Cout_A25_B9;
    full_adder add_a25_b9(P_A25_B9, Cout_A25_B9, P_A26_B8, AND_A25_B9, Cout_A25_B8);

    wire AND_A26_B9;
    and and_a26_b9(AND_A26_B9, A[26], B[9]);
    wire P_A26_B9, Cout_A26_B9;
    full_adder add_a26_b9(P_A26_B9, Cout_A26_B9, P_A27_B8, AND_A26_B9, Cout_A26_B8);

    wire AND_A27_B9;
    and and_a27_b9(AND_A27_B9, A[27], B[9]);
    wire P_A27_B9, Cout_A27_B9;
    full_adder add_a27_b9(P_A27_B9, Cout_A27_B9, P_A28_B8, AND_A27_B9, Cout_A27_B8);

    wire AND_A28_B9;
    and and_a28_b9(AND_A28_B9, A[28], B[9]);
    wire P_A28_B9, Cout_A28_B9;
    full_adder add_a28_b9(P_A28_B9, Cout_A28_B9, P_A29_B8, AND_A28_B9, Cout_A28_B8);

    wire AND_A29_B9;
    and and_a29_b9(AND_A29_B9, A[29], B[9]);
    wire P_A29_B9, Cout_A29_B9;
    full_adder add_a29_b9(P_A29_B9, Cout_A29_B9, P_A30_B8, AND_A29_B9, Cout_A29_B8);

    wire AND_A30_B9;
    and and_a30_b9(AND_A30_B9, A[30], B[9]);
    wire P_A30_B9, Cout_A30_B9;
    full_adder add_a30_b9(P_A30_B9, Cout_A30_B9, P_A31_B8, AND_A30_B9, Cout_A30_B8);

    wire AND_A31_B9;
    nand and_a31_b9(AND_A31_B9, A[31], B[9]);
    wire P_A31_B9, Cout_A31_B9;
    half_adder add_a31_b9(P_A31_B9, Cout_A31_B9, AND_A31_B9, Cout_A31_B8);

    wire AND_A0_B10;
    and and_a0_b10(AND_A0_B10, A[0], B[10]);
    wire P_A0_B10, Cout_A0_B10;
    full_adder add_a0_b10(P_A0_B10, Cout_A0_B10, P_A1_B9, AND_A0_B10, Cout_A0_B9);

    wire AND_A1_B10;
    and and_a1_b10(AND_A1_B10, A[1], B[10]);
    wire P_A1_B10, Cout_A1_B10;
    full_adder add_a1_b10(P_A1_B10, Cout_A1_B10, P_A2_B9, AND_A1_B10, Cout_A1_B9);

    wire AND_A2_B10;
    and and_a2_b10(AND_A2_B10, A[2], B[10]);
    wire P_A2_B10, Cout_A2_B10;
    full_adder add_a2_b10(P_A2_B10, Cout_A2_B10, P_A3_B9, AND_A2_B10, Cout_A2_B9);

    wire AND_A3_B10;
    and and_a3_b10(AND_A3_B10, A[3], B[10]);
    wire P_A3_B10, Cout_A3_B10;
    full_adder add_a3_b10(P_A3_B10, Cout_A3_B10, P_A4_B9, AND_A3_B10, Cout_A3_B9);

    wire AND_A4_B10;
    and and_a4_b10(AND_A4_B10, A[4], B[10]);
    wire P_A4_B10, Cout_A4_B10;
    full_adder add_a4_b10(P_A4_B10, Cout_A4_B10, P_A5_B9, AND_A4_B10, Cout_A4_B9);

    wire AND_A5_B10;
    and and_a5_b10(AND_A5_B10, A[5], B[10]);
    wire P_A5_B10, Cout_A5_B10;
    full_adder add_a5_b10(P_A5_B10, Cout_A5_B10, P_A6_B9, AND_A5_B10, Cout_A5_B9);

    wire AND_A6_B10;
    and and_a6_b10(AND_A6_B10, A[6], B[10]);
    wire P_A6_B10, Cout_A6_B10;
    full_adder add_a6_b10(P_A6_B10, Cout_A6_B10, P_A7_B9, AND_A6_B10, Cout_A6_B9);

    wire AND_A7_B10;
    and and_a7_b10(AND_A7_B10, A[7], B[10]);
    wire P_A7_B10, Cout_A7_B10;
    full_adder add_a7_b10(P_A7_B10, Cout_A7_B10, P_A8_B9, AND_A7_B10, Cout_A7_B9);

    wire AND_A8_B10;
    and and_a8_b10(AND_A8_B10, A[8], B[10]);
    wire P_A8_B10, Cout_A8_B10;
    full_adder add_a8_b10(P_A8_B10, Cout_A8_B10, P_A9_B9, AND_A8_B10, Cout_A8_B9);

    wire AND_A9_B10;
    and and_a9_b10(AND_A9_B10, A[9], B[10]);
    wire P_A9_B10, Cout_A9_B10;
    full_adder add_a9_b10(P_A9_B10, Cout_A9_B10, P_A10_B9, AND_A9_B10, Cout_A9_B9);

    wire AND_A10_B10;
    and and_a10_b10(AND_A10_B10, A[10], B[10]);
    wire P_A10_B10, Cout_A10_B10;
    full_adder add_a10_b10(P_A10_B10, Cout_A10_B10, P_A11_B9, AND_A10_B10, Cout_A10_B9);

    wire AND_A11_B10;
    and and_a11_b10(AND_A11_B10, A[11], B[10]);
    wire P_A11_B10, Cout_A11_B10;
    full_adder add_a11_b10(P_A11_B10, Cout_A11_B10, P_A12_B9, AND_A11_B10, Cout_A11_B9);

    wire AND_A12_B10;
    and and_a12_b10(AND_A12_B10, A[12], B[10]);
    wire P_A12_B10, Cout_A12_B10;
    full_adder add_a12_b10(P_A12_B10, Cout_A12_B10, P_A13_B9, AND_A12_B10, Cout_A12_B9);

    wire AND_A13_B10;
    and and_a13_b10(AND_A13_B10, A[13], B[10]);
    wire P_A13_B10, Cout_A13_B10;
    full_adder add_a13_b10(P_A13_B10, Cout_A13_B10, P_A14_B9, AND_A13_B10, Cout_A13_B9);

    wire AND_A14_B10;
    and and_a14_b10(AND_A14_B10, A[14], B[10]);
    wire P_A14_B10, Cout_A14_B10;
    full_adder add_a14_b10(P_A14_B10, Cout_A14_B10, P_A15_B9, AND_A14_B10, Cout_A14_B9);

    wire AND_A15_B10;
    and and_a15_b10(AND_A15_B10, A[15], B[10]);
    wire P_A15_B10, Cout_A15_B10;
    full_adder add_a15_b10(P_A15_B10, Cout_A15_B10, P_A16_B9, AND_A15_B10, Cout_A15_B9);

    wire AND_A16_B10;
    and and_a16_b10(AND_A16_B10, A[16], B[10]);
    wire P_A16_B10, Cout_A16_B10;
    full_adder add_a16_b10(P_A16_B10, Cout_A16_B10, P_A17_B9, AND_A16_B10, Cout_A16_B9);

    wire AND_A17_B10;
    and and_a17_b10(AND_A17_B10, A[17], B[10]);
    wire P_A17_B10, Cout_A17_B10;
    full_adder add_a17_b10(P_A17_B10, Cout_A17_B10, P_A18_B9, AND_A17_B10, Cout_A17_B9);

    wire AND_A18_B10;
    and and_a18_b10(AND_A18_B10, A[18], B[10]);
    wire P_A18_B10, Cout_A18_B10;
    full_adder add_a18_b10(P_A18_B10, Cout_A18_B10, P_A19_B9, AND_A18_B10, Cout_A18_B9);

    wire AND_A19_B10;
    and and_a19_b10(AND_A19_B10, A[19], B[10]);
    wire P_A19_B10, Cout_A19_B10;
    full_adder add_a19_b10(P_A19_B10, Cout_A19_B10, P_A20_B9, AND_A19_B10, Cout_A19_B9);

    wire AND_A20_B10;
    and and_a20_b10(AND_A20_B10, A[20], B[10]);
    wire P_A20_B10, Cout_A20_B10;
    full_adder add_a20_b10(P_A20_B10, Cout_A20_B10, P_A21_B9, AND_A20_B10, Cout_A20_B9);

    wire AND_A21_B10;
    and and_a21_b10(AND_A21_B10, A[21], B[10]);
    wire P_A21_B10, Cout_A21_B10;
    full_adder add_a21_b10(P_A21_B10, Cout_A21_B10, P_A22_B9, AND_A21_B10, Cout_A21_B9);

    wire AND_A22_B10;
    and and_a22_b10(AND_A22_B10, A[22], B[10]);
    wire P_A22_B10, Cout_A22_B10;
    full_adder add_a22_b10(P_A22_B10, Cout_A22_B10, P_A23_B9, AND_A22_B10, Cout_A22_B9);

    wire AND_A23_B10;
    and and_a23_b10(AND_A23_B10, A[23], B[10]);
    wire P_A23_B10, Cout_A23_B10;
    full_adder add_a23_b10(P_A23_B10, Cout_A23_B10, P_A24_B9, AND_A23_B10, Cout_A23_B9);

    wire AND_A24_B10;
    and and_a24_b10(AND_A24_B10, A[24], B[10]);
    wire P_A24_B10, Cout_A24_B10;
    full_adder add_a24_b10(P_A24_B10, Cout_A24_B10, P_A25_B9, AND_A24_B10, Cout_A24_B9);

    wire AND_A25_B10;
    and and_a25_b10(AND_A25_B10, A[25], B[10]);
    wire P_A25_B10, Cout_A25_B10;
    full_adder add_a25_b10(P_A25_B10, Cout_A25_B10, P_A26_B9, AND_A25_B10, Cout_A25_B9);

    wire AND_A26_B10;
    and and_a26_b10(AND_A26_B10, A[26], B[10]);
    wire P_A26_B10, Cout_A26_B10;
    full_adder add_a26_b10(P_A26_B10, Cout_A26_B10, P_A27_B9, AND_A26_B10, Cout_A26_B9);

    wire AND_A27_B10;
    and and_a27_b10(AND_A27_B10, A[27], B[10]);
    wire P_A27_B10, Cout_A27_B10;
    full_adder add_a27_b10(P_A27_B10, Cout_A27_B10, P_A28_B9, AND_A27_B10, Cout_A27_B9);

    wire AND_A28_B10;
    and and_a28_b10(AND_A28_B10, A[28], B[10]);
    wire P_A28_B10, Cout_A28_B10;
    full_adder add_a28_b10(P_A28_B10, Cout_A28_B10, P_A29_B9, AND_A28_B10, Cout_A28_B9);

    wire AND_A29_B10;
    and and_a29_b10(AND_A29_B10, A[29], B[10]);
    wire P_A29_B10, Cout_A29_B10;
    full_adder add_a29_b10(P_A29_B10, Cout_A29_B10, P_A30_B9, AND_A29_B10, Cout_A29_B9);

    wire AND_A30_B10;
    and and_a30_b10(AND_A30_B10, A[30], B[10]);
    wire P_A30_B10, Cout_A30_B10;
    full_adder add_a30_b10(P_A30_B10, Cout_A30_B10, P_A31_B9, AND_A30_B10, Cout_A30_B9);

    wire AND_A31_B10;
    nand and_a31_b10(AND_A31_B10, A[31], B[10]);
    wire P_A31_B10, Cout_A31_B10;
    half_adder add_a31_b10(P_A31_B10, Cout_A31_B10, AND_A31_B10, Cout_A31_B9);

    wire AND_A0_B11;
    and and_a0_b11(AND_A0_B11, A[0], B[11]);
    wire P_A0_B11, Cout_A0_B11;
    full_adder add_a0_b11(P_A0_B11, Cout_A0_B11, P_A1_B10, AND_A0_B11, Cout_A0_B10);

    wire AND_A1_B11;
    and and_a1_b11(AND_A1_B11, A[1], B[11]);
    wire P_A1_B11, Cout_A1_B11;
    full_adder add_a1_b11(P_A1_B11, Cout_A1_B11, P_A2_B10, AND_A1_B11, Cout_A1_B10);

    wire AND_A2_B11;
    and and_a2_b11(AND_A2_B11, A[2], B[11]);
    wire P_A2_B11, Cout_A2_B11;
    full_adder add_a2_b11(P_A2_B11, Cout_A2_B11, P_A3_B10, AND_A2_B11, Cout_A2_B10);

    wire AND_A3_B11;
    and and_a3_b11(AND_A3_B11, A[3], B[11]);
    wire P_A3_B11, Cout_A3_B11;
    full_adder add_a3_b11(P_A3_B11, Cout_A3_B11, P_A4_B10, AND_A3_B11, Cout_A3_B10);

    wire AND_A4_B11;
    and and_a4_b11(AND_A4_B11, A[4], B[11]);
    wire P_A4_B11, Cout_A4_B11;
    full_adder add_a4_b11(P_A4_B11, Cout_A4_B11, P_A5_B10, AND_A4_B11, Cout_A4_B10);

    wire AND_A5_B11;
    and and_a5_b11(AND_A5_B11, A[5], B[11]);
    wire P_A5_B11, Cout_A5_B11;
    full_adder add_a5_b11(P_A5_B11, Cout_A5_B11, P_A6_B10, AND_A5_B11, Cout_A5_B10);

    wire AND_A6_B11;
    and and_a6_b11(AND_A6_B11, A[6], B[11]);
    wire P_A6_B11, Cout_A6_B11;
    full_adder add_a6_b11(P_A6_B11, Cout_A6_B11, P_A7_B10, AND_A6_B11, Cout_A6_B10);

    wire AND_A7_B11;
    and and_a7_b11(AND_A7_B11, A[7], B[11]);
    wire P_A7_B11, Cout_A7_B11;
    full_adder add_a7_b11(P_A7_B11, Cout_A7_B11, P_A8_B10, AND_A7_B11, Cout_A7_B10);

    wire AND_A8_B11;
    and and_a8_b11(AND_A8_B11, A[8], B[11]);
    wire P_A8_B11, Cout_A8_B11;
    full_adder add_a8_b11(P_A8_B11, Cout_A8_B11, P_A9_B10, AND_A8_B11, Cout_A8_B10);

    wire AND_A9_B11;
    and and_a9_b11(AND_A9_B11, A[9], B[11]);
    wire P_A9_B11, Cout_A9_B11;
    full_adder add_a9_b11(P_A9_B11, Cout_A9_B11, P_A10_B10, AND_A9_B11, Cout_A9_B10);

    wire AND_A10_B11;
    and and_a10_b11(AND_A10_B11, A[10], B[11]);
    wire P_A10_B11, Cout_A10_B11;
    full_adder add_a10_b11(P_A10_B11, Cout_A10_B11, P_A11_B10, AND_A10_B11, Cout_A10_B10);

    wire AND_A11_B11;
    and and_a11_b11(AND_A11_B11, A[11], B[11]);
    wire P_A11_B11, Cout_A11_B11;
    full_adder add_a11_b11(P_A11_B11, Cout_A11_B11, P_A12_B10, AND_A11_B11, Cout_A11_B10);

    wire AND_A12_B11;
    and and_a12_b11(AND_A12_B11, A[12], B[11]);
    wire P_A12_B11, Cout_A12_B11;
    full_adder add_a12_b11(P_A12_B11, Cout_A12_B11, P_A13_B10, AND_A12_B11, Cout_A12_B10);

    wire AND_A13_B11;
    and and_a13_b11(AND_A13_B11, A[13], B[11]);
    wire P_A13_B11, Cout_A13_B11;
    full_adder add_a13_b11(P_A13_B11, Cout_A13_B11, P_A14_B10, AND_A13_B11, Cout_A13_B10);

    wire AND_A14_B11;
    and and_a14_b11(AND_A14_B11, A[14], B[11]);
    wire P_A14_B11, Cout_A14_B11;
    full_adder add_a14_b11(P_A14_B11, Cout_A14_B11, P_A15_B10, AND_A14_B11, Cout_A14_B10);

    wire AND_A15_B11;
    and and_a15_b11(AND_A15_B11, A[15], B[11]);
    wire P_A15_B11, Cout_A15_B11;
    full_adder add_a15_b11(P_A15_B11, Cout_A15_B11, P_A16_B10, AND_A15_B11, Cout_A15_B10);

    wire AND_A16_B11;
    and and_a16_b11(AND_A16_B11, A[16], B[11]);
    wire P_A16_B11, Cout_A16_B11;
    full_adder add_a16_b11(P_A16_B11, Cout_A16_B11, P_A17_B10, AND_A16_B11, Cout_A16_B10);

    wire AND_A17_B11;
    and and_a17_b11(AND_A17_B11, A[17], B[11]);
    wire P_A17_B11, Cout_A17_B11;
    full_adder add_a17_b11(P_A17_B11, Cout_A17_B11, P_A18_B10, AND_A17_B11, Cout_A17_B10);

    wire AND_A18_B11;
    and and_a18_b11(AND_A18_B11, A[18], B[11]);
    wire P_A18_B11, Cout_A18_B11;
    full_adder add_a18_b11(P_A18_B11, Cout_A18_B11, P_A19_B10, AND_A18_B11, Cout_A18_B10);

    wire AND_A19_B11;
    and and_a19_b11(AND_A19_B11, A[19], B[11]);
    wire P_A19_B11, Cout_A19_B11;
    full_adder add_a19_b11(P_A19_B11, Cout_A19_B11, P_A20_B10, AND_A19_B11, Cout_A19_B10);

    wire AND_A20_B11;
    and and_a20_b11(AND_A20_B11, A[20], B[11]);
    wire P_A20_B11, Cout_A20_B11;
    full_adder add_a20_b11(P_A20_B11, Cout_A20_B11, P_A21_B10, AND_A20_B11, Cout_A20_B10);

    wire AND_A21_B11;
    and and_a21_b11(AND_A21_B11, A[21], B[11]);
    wire P_A21_B11, Cout_A21_B11;
    full_adder add_a21_b11(P_A21_B11, Cout_A21_B11, P_A22_B10, AND_A21_B11, Cout_A21_B10);

    wire AND_A22_B11;
    and and_a22_b11(AND_A22_B11, A[22], B[11]);
    wire P_A22_B11, Cout_A22_B11;
    full_adder add_a22_b11(P_A22_B11, Cout_A22_B11, P_A23_B10, AND_A22_B11, Cout_A22_B10);

    wire AND_A23_B11;
    and and_a23_b11(AND_A23_B11, A[23], B[11]);
    wire P_A23_B11, Cout_A23_B11;
    full_adder add_a23_b11(P_A23_B11, Cout_A23_B11, P_A24_B10, AND_A23_B11, Cout_A23_B10);

    wire AND_A24_B11;
    and and_a24_b11(AND_A24_B11, A[24], B[11]);
    wire P_A24_B11, Cout_A24_B11;
    full_adder add_a24_b11(P_A24_B11, Cout_A24_B11, P_A25_B10, AND_A24_B11, Cout_A24_B10);

    wire AND_A25_B11;
    and and_a25_b11(AND_A25_B11, A[25], B[11]);
    wire P_A25_B11, Cout_A25_B11;
    full_adder add_a25_b11(P_A25_B11, Cout_A25_B11, P_A26_B10, AND_A25_B11, Cout_A25_B10);

    wire AND_A26_B11;
    and and_a26_b11(AND_A26_B11, A[26], B[11]);
    wire P_A26_B11, Cout_A26_B11;
    full_adder add_a26_b11(P_A26_B11, Cout_A26_B11, P_A27_B10, AND_A26_B11, Cout_A26_B10);

    wire AND_A27_B11;
    and and_a27_b11(AND_A27_B11, A[27], B[11]);
    wire P_A27_B11, Cout_A27_B11;
    full_adder add_a27_b11(P_A27_B11, Cout_A27_B11, P_A28_B10, AND_A27_B11, Cout_A27_B10);

    wire AND_A28_B11;
    and and_a28_b11(AND_A28_B11, A[28], B[11]);
    wire P_A28_B11, Cout_A28_B11;
    full_adder add_a28_b11(P_A28_B11, Cout_A28_B11, P_A29_B10, AND_A28_B11, Cout_A28_B10);

    wire AND_A29_B11;
    and and_a29_b11(AND_A29_B11, A[29], B[11]);
    wire P_A29_B11, Cout_A29_B11;
    full_adder add_a29_b11(P_A29_B11, Cout_A29_B11, P_A30_B10, AND_A29_B11, Cout_A29_B10);

    wire AND_A30_B11;
    and and_a30_b11(AND_A30_B11, A[30], B[11]);
    wire P_A30_B11, Cout_A30_B11;
    full_adder add_a30_b11(P_A30_B11, Cout_A30_B11, P_A31_B10, AND_A30_B11, Cout_A30_B10);

    wire AND_A31_B11;
    nand and_a31_b11(AND_A31_B11, A[31], B[11]);
    wire P_A31_B11, Cout_A31_B11;
    half_adder add_a31_b11(P_A31_B11, Cout_A31_B11, AND_A31_B11, Cout_A31_B10);

    wire AND_A0_B12;
    and and_a0_b12(AND_A0_B12, A[0], B[12]);
    wire P_A0_B12, Cout_A0_B12;
    full_adder add_a0_b12(P_A0_B12, Cout_A0_B12, P_A1_B11, AND_A0_B12, Cout_A0_B11);

    wire AND_A1_B12;
    and and_a1_b12(AND_A1_B12, A[1], B[12]);
    wire P_A1_B12, Cout_A1_B12;
    full_adder add_a1_b12(P_A1_B12, Cout_A1_B12, P_A2_B11, AND_A1_B12, Cout_A1_B11);

    wire AND_A2_B12;
    and and_a2_b12(AND_A2_B12, A[2], B[12]);
    wire P_A2_B12, Cout_A2_B12;
    full_adder add_a2_b12(P_A2_B12, Cout_A2_B12, P_A3_B11, AND_A2_B12, Cout_A2_B11);

    wire AND_A3_B12;
    and and_a3_b12(AND_A3_B12, A[3], B[12]);
    wire P_A3_B12, Cout_A3_B12;
    full_adder add_a3_b12(P_A3_B12, Cout_A3_B12, P_A4_B11, AND_A3_B12, Cout_A3_B11);

    wire AND_A4_B12;
    and and_a4_b12(AND_A4_B12, A[4], B[12]);
    wire P_A4_B12, Cout_A4_B12;
    full_adder add_a4_b12(P_A4_B12, Cout_A4_B12, P_A5_B11, AND_A4_B12, Cout_A4_B11);

    wire AND_A5_B12;
    and and_a5_b12(AND_A5_B12, A[5], B[12]);
    wire P_A5_B12, Cout_A5_B12;
    full_adder add_a5_b12(P_A5_B12, Cout_A5_B12, P_A6_B11, AND_A5_B12, Cout_A5_B11);

    wire AND_A6_B12;
    and and_a6_b12(AND_A6_B12, A[6], B[12]);
    wire P_A6_B12, Cout_A6_B12;
    full_adder add_a6_b12(P_A6_B12, Cout_A6_B12, P_A7_B11, AND_A6_B12, Cout_A6_B11);

    wire AND_A7_B12;
    and and_a7_b12(AND_A7_B12, A[7], B[12]);
    wire P_A7_B12, Cout_A7_B12;
    full_adder add_a7_b12(P_A7_B12, Cout_A7_B12, P_A8_B11, AND_A7_B12, Cout_A7_B11);

    wire AND_A8_B12;
    and and_a8_b12(AND_A8_B12, A[8], B[12]);
    wire P_A8_B12, Cout_A8_B12;
    full_adder add_a8_b12(P_A8_B12, Cout_A8_B12, P_A9_B11, AND_A8_B12, Cout_A8_B11);

    wire AND_A9_B12;
    and and_a9_b12(AND_A9_B12, A[9], B[12]);
    wire P_A9_B12, Cout_A9_B12;
    full_adder add_a9_b12(P_A9_B12, Cout_A9_B12, P_A10_B11, AND_A9_B12, Cout_A9_B11);

    wire AND_A10_B12;
    and and_a10_b12(AND_A10_B12, A[10], B[12]);
    wire P_A10_B12, Cout_A10_B12;
    full_adder add_a10_b12(P_A10_B12, Cout_A10_B12, P_A11_B11, AND_A10_B12, Cout_A10_B11);

    wire AND_A11_B12;
    and and_a11_b12(AND_A11_B12, A[11], B[12]);
    wire P_A11_B12, Cout_A11_B12;
    full_adder add_a11_b12(P_A11_B12, Cout_A11_B12, P_A12_B11, AND_A11_B12, Cout_A11_B11);

    wire AND_A12_B12;
    and and_a12_b12(AND_A12_B12, A[12], B[12]);
    wire P_A12_B12, Cout_A12_B12;
    full_adder add_a12_b12(P_A12_B12, Cout_A12_B12, P_A13_B11, AND_A12_B12, Cout_A12_B11);

    wire AND_A13_B12;
    and and_a13_b12(AND_A13_B12, A[13], B[12]);
    wire P_A13_B12, Cout_A13_B12;
    full_adder add_a13_b12(P_A13_B12, Cout_A13_B12, P_A14_B11, AND_A13_B12, Cout_A13_B11);

    wire AND_A14_B12;
    and and_a14_b12(AND_A14_B12, A[14], B[12]);
    wire P_A14_B12, Cout_A14_B12;
    full_adder add_a14_b12(P_A14_B12, Cout_A14_B12, P_A15_B11, AND_A14_B12, Cout_A14_B11);

    wire AND_A15_B12;
    and and_a15_b12(AND_A15_B12, A[15], B[12]);
    wire P_A15_B12, Cout_A15_B12;
    full_adder add_a15_b12(P_A15_B12, Cout_A15_B12, P_A16_B11, AND_A15_B12, Cout_A15_B11);

    wire AND_A16_B12;
    and and_a16_b12(AND_A16_B12, A[16], B[12]);
    wire P_A16_B12, Cout_A16_B12;
    full_adder add_a16_b12(P_A16_B12, Cout_A16_B12, P_A17_B11, AND_A16_B12, Cout_A16_B11);

    wire AND_A17_B12;
    and and_a17_b12(AND_A17_B12, A[17], B[12]);
    wire P_A17_B12, Cout_A17_B12;
    full_adder add_a17_b12(P_A17_B12, Cout_A17_B12, P_A18_B11, AND_A17_B12, Cout_A17_B11);

    wire AND_A18_B12;
    and and_a18_b12(AND_A18_B12, A[18], B[12]);
    wire P_A18_B12, Cout_A18_B12;
    full_adder add_a18_b12(P_A18_B12, Cout_A18_B12, P_A19_B11, AND_A18_B12, Cout_A18_B11);

    wire AND_A19_B12;
    and and_a19_b12(AND_A19_B12, A[19], B[12]);
    wire P_A19_B12, Cout_A19_B12;
    full_adder add_a19_b12(P_A19_B12, Cout_A19_B12, P_A20_B11, AND_A19_B12, Cout_A19_B11);

    wire AND_A20_B12;
    and and_a20_b12(AND_A20_B12, A[20], B[12]);
    wire P_A20_B12, Cout_A20_B12;
    full_adder add_a20_b12(P_A20_B12, Cout_A20_B12, P_A21_B11, AND_A20_B12, Cout_A20_B11);

    wire AND_A21_B12;
    and and_a21_b12(AND_A21_B12, A[21], B[12]);
    wire P_A21_B12, Cout_A21_B12;
    full_adder add_a21_b12(P_A21_B12, Cout_A21_B12, P_A22_B11, AND_A21_B12, Cout_A21_B11);

    wire AND_A22_B12;
    and and_a22_b12(AND_A22_B12, A[22], B[12]);
    wire P_A22_B12, Cout_A22_B12;
    full_adder add_a22_b12(P_A22_B12, Cout_A22_B12, P_A23_B11, AND_A22_B12, Cout_A22_B11);

    wire AND_A23_B12;
    and and_a23_b12(AND_A23_B12, A[23], B[12]);
    wire P_A23_B12, Cout_A23_B12;
    full_adder add_a23_b12(P_A23_B12, Cout_A23_B12, P_A24_B11, AND_A23_B12, Cout_A23_B11);

    wire AND_A24_B12;
    and and_a24_b12(AND_A24_B12, A[24], B[12]);
    wire P_A24_B12, Cout_A24_B12;
    full_adder add_a24_b12(P_A24_B12, Cout_A24_B12, P_A25_B11, AND_A24_B12, Cout_A24_B11);

    wire AND_A25_B12;
    and and_a25_b12(AND_A25_B12, A[25], B[12]);
    wire P_A25_B12, Cout_A25_B12;
    full_adder add_a25_b12(P_A25_B12, Cout_A25_B12, P_A26_B11, AND_A25_B12, Cout_A25_B11);

    wire AND_A26_B12;
    and and_a26_b12(AND_A26_B12, A[26], B[12]);
    wire P_A26_B12, Cout_A26_B12;
    full_adder add_a26_b12(P_A26_B12, Cout_A26_B12, P_A27_B11, AND_A26_B12, Cout_A26_B11);

    wire AND_A27_B12;
    and and_a27_b12(AND_A27_B12, A[27], B[12]);
    wire P_A27_B12, Cout_A27_B12;
    full_adder add_a27_b12(P_A27_B12, Cout_A27_B12, P_A28_B11, AND_A27_B12, Cout_A27_B11);

    wire AND_A28_B12;
    and and_a28_b12(AND_A28_B12, A[28], B[12]);
    wire P_A28_B12, Cout_A28_B12;
    full_adder add_a28_b12(P_A28_B12, Cout_A28_B12, P_A29_B11, AND_A28_B12, Cout_A28_B11);

    wire AND_A29_B12;
    and and_a29_b12(AND_A29_B12, A[29], B[12]);
    wire P_A29_B12, Cout_A29_B12;
    full_adder add_a29_b12(P_A29_B12, Cout_A29_B12, P_A30_B11, AND_A29_B12, Cout_A29_B11);

    wire AND_A30_B12;
    and and_a30_b12(AND_A30_B12, A[30], B[12]);
    wire P_A30_B12, Cout_A30_B12;
    full_adder add_a30_b12(P_A30_B12, Cout_A30_B12, P_A31_B11, AND_A30_B12, Cout_A30_B11);

    wire AND_A31_B12;
    nand and_a31_b12(AND_A31_B12, A[31], B[12]);
    wire P_A31_B12, Cout_A31_B12;
    half_adder add_a31_b12(P_A31_B12, Cout_A31_B12, AND_A31_B12, Cout_A31_B11);

    wire AND_A0_B13;
    and and_a0_b13(AND_A0_B13, A[0], B[13]);
    wire P_A0_B13, Cout_A0_B13;
    full_adder add_a0_b13(P_A0_B13, Cout_A0_B13, P_A1_B12, AND_A0_B13, Cout_A0_B12);

    wire AND_A1_B13;
    and and_a1_b13(AND_A1_B13, A[1], B[13]);
    wire P_A1_B13, Cout_A1_B13;
    full_adder add_a1_b13(P_A1_B13, Cout_A1_B13, P_A2_B12, AND_A1_B13, Cout_A1_B12);

    wire AND_A2_B13;
    and and_a2_b13(AND_A2_B13, A[2], B[13]);
    wire P_A2_B13, Cout_A2_B13;
    full_adder add_a2_b13(P_A2_B13, Cout_A2_B13, P_A3_B12, AND_A2_B13, Cout_A2_B12);

    wire AND_A3_B13;
    and and_a3_b13(AND_A3_B13, A[3], B[13]);
    wire P_A3_B13, Cout_A3_B13;
    full_adder add_a3_b13(P_A3_B13, Cout_A3_B13, P_A4_B12, AND_A3_B13, Cout_A3_B12);

    wire AND_A4_B13;
    and and_a4_b13(AND_A4_B13, A[4], B[13]);
    wire P_A4_B13, Cout_A4_B13;
    full_adder add_a4_b13(P_A4_B13, Cout_A4_B13, P_A5_B12, AND_A4_B13, Cout_A4_B12);

    wire AND_A5_B13;
    and and_a5_b13(AND_A5_B13, A[5], B[13]);
    wire P_A5_B13, Cout_A5_B13;
    full_adder add_a5_b13(P_A5_B13, Cout_A5_B13, P_A6_B12, AND_A5_B13, Cout_A5_B12);

    wire AND_A6_B13;
    and and_a6_b13(AND_A6_B13, A[6], B[13]);
    wire P_A6_B13, Cout_A6_B13;
    full_adder add_a6_b13(P_A6_B13, Cout_A6_B13, P_A7_B12, AND_A6_B13, Cout_A6_B12);

    wire AND_A7_B13;
    and and_a7_b13(AND_A7_B13, A[7], B[13]);
    wire P_A7_B13, Cout_A7_B13;
    full_adder add_a7_b13(P_A7_B13, Cout_A7_B13, P_A8_B12, AND_A7_B13, Cout_A7_B12);

    wire AND_A8_B13;
    and and_a8_b13(AND_A8_B13, A[8], B[13]);
    wire P_A8_B13, Cout_A8_B13;
    full_adder add_a8_b13(P_A8_B13, Cout_A8_B13, P_A9_B12, AND_A8_B13, Cout_A8_B12);

    wire AND_A9_B13;
    and and_a9_b13(AND_A9_B13, A[9], B[13]);
    wire P_A9_B13, Cout_A9_B13;
    full_adder add_a9_b13(P_A9_B13, Cout_A9_B13, P_A10_B12, AND_A9_B13, Cout_A9_B12);

    wire AND_A10_B13;
    and and_a10_b13(AND_A10_B13, A[10], B[13]);
    wire P_A10_B13, Cout_A10_B13;
    full_adder add_a10_b13(P_A10_B13, Cout_A10_B13, P_A11_B12, AND_A10_B13, Cout_A10_B12);

    wire AND_A11_B13;
    and and_a11_b13(AND_A11_B13, A[11], B[13]);
    wire P_A11_B13, Cout_A11_B13;
    full_adder add_a11_b13(P_A11_B13, Cout_A11_B13, P_A12_B12, AND_A11_B13, Cout_A11_B12);

    wire AND_A12_B13;
    and and_a12_b13(AND_A12_B13, A[12], B[13]);
    wire P_A12_B13, Cout_A12_B13;
    full_adder add_a12_b13(P_A12_B13, Cout_A12_B13, P_A13_B12, AND_A12_B13, Cout_A12_B12);

    wire AND_A13_B13;
    and and_a13_b13(AND_A13_B13, A[13], B[13]);
    wire P_A13_B13, Cout_A13_B13;
    full_adder add_a13_b13(P_A13_B13, Cout_A13_B13, P_A14_B12, AND_A13_B13, Cout_A13_B12);

    wire AND_A14_B13;
    and and_a14_b13(AND_A14_B13, A[14], B[13]);
    wire P_A14_B13, Cout_A14_B13;
    full_adder add_a14_b13(P_A14_B13, Cout_A14_B13, P_A15_B12, AND_A14_B13, Cout_A14_B12);

    wire AND_A15_B13;
    and and_a15_b13(AND_A15_B13, A[15], B[13]);
    wire P_A15_B13, Cout_A15_B13;
    full_adder add_a15_b13(P_A15_B13, Cout_A15_B13, P_A16_B12, AND_A15_B13, Cout_A15_B12);

    wire AND_A16_B13;
    and and_a16_b13(AND_A16_B13, A[16], B[13]);
    wire P_A16_B13, Cout_A16_B13;
    full_adder add_a16_b13(P_A16_B13, Cout_A16_B13, P_A17_B12, AND_A16_B13, Cout_A16_B12);

    wire AND_A17_B13;
    and and_a17_b13(AND_A17_B13, A[17], B[13]);
    wire P_A17_B13, Cout_A17_B13;
    full_adder add_a17_b13(P_A17_B13, Cout_A17_B13, P_A18_B12, AND_A17_B13, Cout_A17_B12);

    wire AND_A18_B13;
    and and_a18_b13(AND_A18_B13, A[18], B[13]);
    wire P_A18_B13, Cout_A18_B13;
    full_adder add_a18_b13(P_A18_B13, Cout_A18_B13, P_A19_B12, AND_A18_B13, Cout_A18_B12);

    wire AND_A19_B13;
    and and_a19_b13(AND_A19_B13, A[19], B[13]);
    wire P_A19_B13, Cout_A19_B13;
    full_adder add_a19_b13(P_A19_B13, Cout_A19_B13, P_A20_B12, AND_A19_B13, Cout_A19_B12);

    wire AND_A20_B13;
    and and_a20_b13(AND_A20_B13, A[20], B[13]);
    wire P_A20_B13, Cout_A20_B13;
    full_adder add_a20_b13(P_A20_B13, Cout_A20_B13, P_A21_B12, AND_A20_B13, Cout_A20_B12);

    wire AND_A21_B13;
    and and_a21_b13(AND_A21_B13, A[21], B[13]);
    wire P_A21_B13, Cout_A21_B13;
    full_adder add_a21_b13(P_A21_B13, Cout_A21_B13, P_A22_B12, AND_A21_B13, Cout_A21_B12);

    wire AND_A22_B13;
    and and_a22_b13(AND_A22_B13, A[22], B[13]);
    wire P_A22_B13, Cout_A22_B13;
    full_adder add_a22_b13(P_A22_B13, Cout_A22_B13, P_A23_B12, AND_A22_B13, Cout_A22_B12);

    wire AND_A23_B13;
    and and_a23_b13(AND_A23_B13, A[23], B[13]);
    wire P_A23_B13, Cout_A23_B13;
    full_adder add_a23_b13(P_A23_B13, Cout_A23_B13, P_A24_B12, AND_A23_B13, Cout_A23_B12);

    wire AND_A24_B13;
    and and_a24_b13(AND_A24_B13, A[24], B[13]);
    wire P_A24_B13, Cout_A24_B13;
    full_adder add_a24_b13(P_A24_B13, Cout_A24_B13, P_A25_B12, AND_A24_B13, Cout_A24_B12);

    wire AND_A25_B13;
    and and_a25_b13(AND_A25_B13, A[25], B[13]);
    wire P_A25_B13, Cout_A25_B13;
    full_adder add_a25_b13(P_A25_B13, Cout_A25_B13, P_A26_B12, AND_A25_B13, Cout_A25_B12);

    wire AND_A26_B13;
    and and_a26_b13(AND_A26_B13, A[26], B[13]);
    wire P_A26_B13, Cout_A26_B13;
    full_adder add_a26_b13(P_A26_B13, Cout_A26_B13, P_A27_B12, AND_A26_B13, Cout_A26_B12);

    wire AND_A27_B13;
    and and_a27_b13(AND_A27_B13, A[27], B[13]);
    wire P_A27_B13, Cout_A27_B13;
    full_adder add_a27_b13(P_A27_B13, Cout_A27_B13, P_A28_B12, AND_A27_B13, Cout_A27_B12);

    wire AND_A28_B13;
    and and_a28_b13(AND_A28_B13, A[28], B[13]);
    wire P_A28_B13, Cout_A28_B13;
    full_adder add_a28_b13(P_A28_B13, Cout_A28_B13, P_A29_B12, AND_A28_B13, Cout_A28_B12);

    wire AND_A29_B13;
    and and_a29_b13(AND_A29_B13, A[29], B[13]);
    wire P_A29_B13, Cout_A29_B13;
    full_adder add_a29_b13(P_A29_B13, Cout_A29_B13, P_A30_B12, AND_A29_B13, Cout_A29_B12);

    wire AND_A30_B13;
    and and_a30_b13(AND_A30_B13, A[30], B[13]);
    wire P_A30_B13, Cout_A30_B13;
    full_adder add_a30_b13(P_A30_B13, Cout_A30_B13, P_A31_B12, AND_A30_B13, Cout_A30_B12);

    wire AND_A31_B13;
    nand and_a31_b13(AND_A31_B13, A[31], B[13]);
    wire P_A31_B13, Cout_A31_B13;
    half_adder add_a31_b13(P_A31_B13, Cout_A31_B13, AND_A31_B13, Cout_A31_B12);

    wire AND_A0_B14;
    and and_a0_b14(AND_A0_B14, A[0], B[14]);
    wire P_A0_B14, Cout_A0_B14;
    full_adder add_a0_b14(P_A0_B14, Cout_A0_B14, P_A1_B13, AND_A0_B14, Cout_A0_B13);

    wire AND_A1_B14;
    and and_a1_b14(AND_A1_B14, A[1], B[14]);
    wire P_A1_B14, Cout_A1_B14;
    full_adder add_a1_b14(P_A1_B14, Cout_A1_B14, P_A2_B13, AND_A1_B14, Cout_A1_B13);

    wire AND_A2_B14;
    and and_a2_b14(AND_A2_B14, A[2], B[14]);
    wire P_A2_B14, Cout_A2_B14;
    full_adder add_a2_b14(P_A2_B14, Cout_A2_B14, P_A3_B13, AND_A2_B14, Cout_A2_B13);

    wire AND_A3_B14;
    and and_a3_b14(AND_A3_B14, A[3], B[14]);
    wire P_A3_B14, Cout_A3_B14;
    full_adder add_a3_b14(P_A3_B14, Cout_A3_B14, P_A4_B13, AND_A3_B14, Cout_A3_B13);

    wire AND_A4_B14;
    and and_a4_b14(AND_A4_B14, A[4], B[14]);
    wire P_A4_B14, Cout_A4_B14;
    full_adder add_a4_b14(P_A4_B14, Cout_A4_B14, P_A5_B13, AND_A4_B14, Cout_A4_B13);

    wire AND_A5_B14;
    and and_a5_b14(AND_A5_B14, A[5], B[14]);
    wire P_A5_B14, Cout_A5_B14;
    full_adder add_a5_b14(P_A5_B14, Cout_A5_B14, P_A6_B13, AND_A5_B14, Cout_A5_B13);

    wire AND_A6_B14;
    and and_a6_b14(AND_A6_B14, A[6], B[14]);
    wire P_A6_B14, Cout_A6_B14;
    full_adder add_a6_b14(P_A6_B14, Cout_A6_B14, P_A7_B13, AND_A6_B14, Cout_A6_B13);

    wire AND_A7_B14;
    and and_a7_b14(AND_A7_B14, A[7], B[14]);
    wire P_A7_B14, Cout_A7_B14;
    full_adder add_a7_b14(P_A7_B14, Cout_A7_B14, P_A8_B13, AND_A7_B14, Cout_A7_B13);

    wire AND_A8_B14;
    and and_a8_b14(AND_A8_B14, A[8], B[14]);
    wire P_A8_B14, Cout_A8_B14;
    full_adder add_a8_b14(P_A8_B14, Cout_A8_B14, P_A9_B13, AND_A8_B14, Cout_A8_B13);

    wire AND_A9_B14;
    and and_a9_b14(AND_A9_B14, A[9], B[14]);
    wire P_A9_B14, Cout_A9_B14;
    full_adder add_a9_b14(P_A9_B14, Cout_A9_B14, P_A10_B13, AND_A9_B14, Cout_A9_B13);

    wire AND_A10_B14;
    and and_a10_b14(AND_A10_B14, A[10], B[14]);
    wire P_A10_B14, Cout_A10_B14;
    full_adder add_a10_b14(P_A10_B14, Cout_A10_B14, P_A11_B13, AND_A10_B14, Cout_A10_B13);

    wire AND_A11_B14;
    and and_a11_b14(AND_A11_B14, A[11], B[14]);
    wire P_A11_B14, Cout_A11_B14;
    full_adder add_a11_b14(P_A11_B14, Cout_A11_B14, P_A12_B13, AND_A11_B14, Cout_A11_B13);

    wire AND_A12_B14;
    and and_a12_b14(AND_A12_B14, A[12], B[14]);
    wire P_A12_B14, Cout_A12_B14;
    full_adder add_a12_b14(P_A12_B14, Cout_A12_B14, P_A13_B13, AND_A12_B14, Cout_A12_B13);

    wire AND_A13_B14;
    and and_a13_b14(AND_A13_B14, A[13], B[14]);
    wire P_A13_B14, Cout_A13_B14;
    full_adder add_a13_b14(P_A13_B14, Cout_A13_B14, P_A14_B13, AND_A13_B14, Cout_A13_B13);

    wire AND_A14_B14;
    and and_a14_b14(AND_A14_B14, A[14], B[14]);
    wire P_A14_B14, Cout_A14_B14;
    full_adder add_a14_b14(P_A14_B14, Cout_A14_B14, P_A15_B13, AND_A14_B14, Cout_A14_B13);

    wire AND_A15_B14;
    and and_a15_b14(AND_A15_B14, A[15], B[14]);
    wire P_A15_B14, Cout_A15_B14;
    full_adder add_a15_b14(P_A15_B14, Cout_A15_B14, P_A16_B13, AND_A15_B14, Cout_A15_B13);

    wire AND_A16_B14;
    and and_a16_b14(AND_A16_B14, A[16], B[14]);
    wire P_A16_B14, Cout_A16_B14;
    full_adder add_a16_b14(P_A16_B14, Cout_A16_B14, P_A17_B13, AND_A16_B14, Cout_A16_B13);

    wire AND_A17_B14;
    and and_a17_b14(AND_A17_B14, A[17], B[14]);
    wire P_A17_B14, Cout_A17_B14;
    full_adder add_a17_b14(P_A17_B14, Cout_A17_B14, P_A18_B13, AND_A17_B14, Cout_A17_B13);

    wire AND_A18_B14;
    and and_a18_b14(AND_A18_B14, A[18], B[14]);
    wire P_A18_B14, Cout_A18_B14;
    full_adder add_a18_b14(P_A18_B14, Cout_A18_B14, P_A19_B13, AND_A18_B14, Cout_A18_B13);

    wire AND_A19_B14;
    and and_a19_b14(AND_A19_B14, A[19], B[14]);
    wire P_A19_B14, Cout_A19_B14;
    full_adder add_a19_b14(P_A19_B14, Cout_A19_B14, P_A20_B13, AND_A19_B14, Cout_A19_B13);

    wire AND_A20_B14;
    and and_a20_b14(AND_A20_B14, A[20], B[14]);
    wire P_A20_B14, Cout_A20_B14;
    full_adder add_a20_b14(P_A20_B14, Cout_A20_B14, P_A21_B13, AND_A20_B14, Cout_A20_B13);

    wire AND_A21_B14;
    and and_a21_b14(AND_A21_B14, A[21], B[14]);
    wire P_A21_B14, Cout_A21_B14;
    full_adder add_a21_b14(P_A21_B14, Cout_A21_B14, P_A22_B13, AND_A21_B14, Cout_A21_B13);

    wire AND_A22_B14;
    and and_a22_b14(AND_A22_B14, A[22], B[14]);
    wire P_A22_B14, Cout_A22_B14;
    full_adder add_a22_b14(P_A22_B14, Cout_A22_B14, P_A23_B13, AND_A22_B14, Cout_A22_B13);

    wire AND_A23_B14;
    and and_a23_b14(AND_A23_B14, A[23], B[14]);
    wire P_A23_B14, Cout_A23_B14;
    full_adder add_a23_b14(P_A23_B14, Cout_A23_B14, P_A24_B13, AND_A23_B14, Cout_A23_B13);

    wire AND_A24_B14;
    and and_a24_b14(AND_A24_B14, A[24], B[14]);
    wire P_A24_B14, Cout_A24_B14;
    full_adder add_a24_b14(P_A24_B14, Cout_A24_B14, P_A25_B13, AND_A24_B14, Cout_A24_B13);

    wire AND_A25_B14;
    and and_a25_b14(AND_A25_B14, A[25], B[14]);
    wire P_A25_B14, Cout_A25_B14;
    full_adder add_a25_b14(P_A25_B14, Cout_A25_B14, P_A26_B13, AND_A25_B14, Cout_A25_B13);

    wire AND_A26_B14;
    and and_a26_b14(AND_A26_B14, A[26], B[14]);
    wire P_A26_B14, Cout_A26_B14;
    full_adder add_a26_b14(P_A26_B14, Cout_A26_B14, P_A27_B13, AND_A26_B14, Cout_A26_B13);

    wire AND_A27_B14;
    and and_a27_b14(AND_A27_B14, A[27], B[14]);
    wire P_A27_B14, Cout_A27_B14;
    full_adder add_a27_b14(P_A27_B14, Cout_A27_B14, P_A28_B13, AND_A27_B14, Cout_A27_B13);

    wire AND_A28_B14;
    and and_a28_b14(AND_A28_B14, A[28], B[14]);
    wire P_A28_B14, Cout_A28_B14;
    full_adder add_a28_b14(P_A28_B14, Cout_A28_B14, P_A29_B13, AND_A28_B14, Cout_A28_B13);

    wire AND_A29_B14;
    and and_a29_b14(AND_A29_B14, A[29], B[14]);
    wire P_A29_B14, Cout_A29_B14;
    full_adder add_a29_b14(P_A29_B14, Cout_A29_B14, P_A30_B13, AND_A29_B14, Cout_A29_B13);

    wire AND_A30_B14;
    and and_a30_b14(AND_A30_B14, A[30], B[14]);
    wire P_A30_B14, Cout_A30_B14;
    full_adder add_a30_b14(P_A30_B14, Cout_A30_B14, P_A31_B13, AND_A30_B14, Cout_A30_B13);

    wire AND_A31_B14;
    nand and_a31_b14(AND_A31_B14, A[31], B[14]);
    wire P_A31_B14, Cout_A31_B14;
    half_adder add_a31_b14(P_A31_B14, Cout_A31_B14, AND_A31_B14, Cout_A31_B13);

    wire AND_A0_B15;
    and and_a0_b15(AND_A0_B15, A[0], B[15]);
    wire P_A0_B15, Cout_A0_B15;
    full_adder add_a0_b15(P_A0_B15, Cout_A0_B15, P_A1_B14, AND_A0_B15, Cout_A0_B14);

    wire AND_A1_B15;
    and and_a1_b15(AND_A1_B15, A[1], B[15]);
    wire P_A1_B15, Cout_A1_B15;
    full_adder add_a1_b15(P_A1_B15, Cout_A1_B15, P_A2_B14, AND_A1_B15, Cout_A1_B14);

    wire AND_A2_B15;
    and and_a2_b15(AND_A2_B15, A[2], B[15]);
    wire P_A2_B15, Cout_A2_B15;
    full_adder add_a2_b15(P_A2_B15, Cout_A2_B15, P_A3_B14, AND_A2_B15, Cout_A2_B14);

    wire AND_A3_B15;
    and and_a3_b15(AND_A3_B15, A[3], B[15]);
    wire P_A3_B15, Cout_A3_B15;
    full_adder add_a3_b15(P_A3_B15, Cout_A3_B15, P_A4_B14, AND_A3_B15, Cout_A3_B14);

    wire AND_A4_B15;
    and and_a4_b15(AND_A4_B15, A[4], B[15]);
    wire P_A4_B15, Cout_A4_B15;
    full_adder add_a4_b15(P_A4_B15, Cout_A4_B15, P_A5_B14, AND_A4_B15, Cout_A4_B14);

    wire AND_A5_B15;
    and and_a5_b15(AND_A5_B15, A[5], B[15]);
    wire P_A5_B15, Cout_A5_B15;
    full_adder add_a5_b15(P_A5_B15, Cout_A5_B15, P_A6_B14, AND_A5_B15, Cout_A5_B14);

    wire AND_A6_B15;
    and and_a6_b15(AND_A6_B15, A[6], B[15]);
    wire P_A6_B15, Cout_A6_B15;
    full_adder add_a6_b15(P_A6_B15, Cout_A6_B15, P_A7_B14, AND_A6_B15, Cout_A6_B14);

    wire AND_A7_B15;
    and and_a7_b15(AND_A7_B15, A[7], B[15]);
    wire P_A7_B15, Cout_A7_B15;
    full_adder add_a7_b15(P_A7_B15, Cout_A7_B15, P_A8_B14, AND_A7_B15, Cout_A7_B14);

    wire AND_A8_B15;
    and and_a8_b15(AND_A8_B15, A[8], B[15]);
    wire P_A8_B15, Cout_A8_B15;
    full_adder add_a8_b15(P_A8_B15, Cout_A8_B15, P_A9_B14, AND_A8_B15, Cout_A8_B14);

    wire AND_A9_B15;
    and and_a9_b15(AND_A9_B15, A[9], B[15]);
    wire P_A9_B15, Cout_A9_B15;
    full_adder add_a9_b15(P_A9_B15, Cout_A9_B15, P_A10_B14, AND_A9_B15, Cout_A9_B14);

    wire AND_A10_B15;
    and and_a10_b15(AND_A10_B15, A[10], B[15]);
    wire P_A10_B15, Cout_A10_B15;
    full_adder add_a10_b15(P_A10_B15, Cout_A10_B15, P_A11_B14, AND_A10_B15, Cout_A10_B14);

    wire AND_A11_B15;
    and and_a11_b15(AND_A11_B15, A[11], B[15]);
    wire P_A11_B15, Cout_A11_B15;
    full_adder add_a11_b15(P_A11_B15, Cout_A11_B15, P_A12_B14, AND_A11_B15, Cout_A11_B14);

    wire AND_A12_B15;
    and and_a12_b15(AND_A12_B15, A[12], B[15]);
    wire P_A12_B15, Cout_A12_B15;
    full_adder add_a12_b15(P_A12_B15, Cout_A12_B15, P_A13_B14, AND_A12_B15, Cout_A12_B14);

    wire AND_A13_B15;
    and and_a13_b15(AND_A13_B15, A[13], B[15]);
    wire P_A13_B15, Cout_A13_B15;
    full_adder add_a13_b15(P_A13_B15, Cout_A13_B15, P_A14_B14, AND_A13_B15, Cout_A13_B14);

    wire AND_A14_B15;
    and and_a14_b15(AND_A14_B15, A[14], B[15]);
    wire P_A14_B15, Cout_A14_B15;
    full_adder add_a14_b15(P_A14_B15, Cout_A14_B15, P_A15_B14, AND_A14_B15, Cout_A14_B14);

    wire AND_A15_B15;
    and and_a15_b15(AND_A15_B15, A[15], B[15]);
    wire P_A15_B15, Cout_A15_B15;
    full_adder add_a15_b15(P_A15_B15, Cout_A15_B15, P_A16_B14, AND_A15_B15, Cout_A15_B14);

    wire AND_A16_B15;
    and and_a16_b15(AND_A16_B15, A[16], B[15]);
    wire P_A16_B15, Cout_A16_B15;
    full_adder add_a16_b15(P_A16_B15, Cout_A16_B15, P_A17_B14, AND_A16_B15, Cout_A16_B14);

    wire AND_A17_B15;
    and and_a17_b15(AND_A17_B15, A[17], B[15]);
    wire P_A17_B15, Cout_A17_B15;
    full_adder add_a17_b15(P_A17_B15, Cout_A17_B15, P_A18_B14, AND_A17_B15, Cout_A17_B14);

    wire AND_A18_B15;
    and and_a18_b15(AND_A18_B15, A[18], B[15]);
    wire P_A18_B15, Cout_A18_B15;
    full_adder add_a18_b15(P_A18_B15, Cout_A18_B15, P_A19_B14, AND_A18_B15, Cout_A18_B14);

    wire AND_A19_B15;
    and and_a19_b15(AND_A19_B15, A[19], B[15]);
    wire P_A19_B15, Cout_A19_B15;
    full_adder add_a19_b15(P_A19_B15, Cout_A19_B15, P_A20_B14, AND_A19_B15, Cout_A19_B14);

    wire AND_A20_B15;
    and and_a20_b15(AND_A20_B15, A[20], B[15]);
    wire P_A20_B15, Cout_A20_B15;
    full_adder add_a20_b15(P_A20_B15, Cout_A20_B15, P_A21_B14, AND_A20_B15, Cout_A20_B14);

    wire AND_A21_B15;
    and and_a21_b15(AND_A21_B15, A[21], B[15]);
    wire P_A21_B15, Cout_A21_B15;
    full_adder add_a21_b15(P_A21_B15, Cout_A21_B15, P_A22_B14, AND_A21_B15, Cout_A21_B14);

    wire AND_A22_B15;
    and and_a22_b15(AND_A22_B15, A[22], B[15]);
    wire P_A22_B15, Cout_A22_B15;
    full_adder add_a22_b15(P_A22_B15, Cout_A22_B15, P_A23_B14, AND_A22_B15, Cout_A22_B14);

    wire AND_A23_B15;
    and and_a23_b15(AND_A23_B15, A[23], B[15]);
    wire P_A23_B15, Cout_A23_B15;
    full_adder add_a23_b15(P_A23_B15, Cout_A23_B15, P_A24_B14, AND_A23_B15, Cout_A23_B14);

    wire AND_A24_B15;
    and and_a24_b15(AND_A24_B15, A[24], B[15]);
    wire P_A24_B15, Cout_A24_B15;
    full_adder add_a24_b15(P_A24_B15, Cout_A24_B15, P_A25_B14, AND_A24_B15, Cout_A24_B14);

    wire AND_A25_B15;
    and and_a25_b15(AND_A25_B15, A[25], B[15]);
    wire P_A25_B15, Cout_A25_B15;
    full_adder add_a25_b15(P_A25_B15, Cout_A25_B15, P_A26_B14, AND_A25_B15, Cout_A25_B14);

    wire AND_A26_B15;
    and and_a26_b15(AND_A26_B15, A[26], B[15]);
    wire P_A26_B15, Cout_A26_B15;
    full_adder add_a26_b15(P_A26_B15, Cout_A26_B15, P_A27_B14, AND_A26_B15, Cout_A26_B14);

    wire AND_A27_B15;
    and and_a27_b15(AND_A27_B15, A[27], B[15]);
    wire P_A27_B15, Cout_A27_B15;
    full_adder add_a27_b15(P_A27_B15, Cout_A27_B15, P_A28_B14, AND_A27_B15, Cout_A27_B14);

    wire AND_A28_B15;
    and and_a28_b15(AND_A28_B15, A[28], B[15]);
    wire P_A28_B15, Cout_A28_B15;
    full_adder add_a28_b15(P_A28_B15, Cout_A28_B15, P_A29_B14, AND_A28_B15, Cout_A28_B14);

    wire AND_A29_B15;
    and and_a29_b15(AND_A29_B15, A[29], B[15]);
    wire P_A29_B15, Cout_A29_B15;
    full_adder add_a29_b15(P_A29_B15, Cout_A29_B15, P_A30_B14, AND_A29_B15, Cout_A29_B14);

    wire AND_A30_B15;
    and and_a30_b15(AND_A30_B15, A[30], B[15]);
    wire P_A30_B15, Cout_A30_B15;
    full_adder add_a30_b15(P_A30_B15, Cout_A30_B15, P_A31_B14, AND_A30_B15, Cout_A30_B14);

    wire AND_A31_B15;
    nand and_a31_b15(AND_A31_B15, A[31], B[15]);
    wire P_A31_B15, Cout_A31_B15;
    half_adder add_a31_b15(P_A31_B15, Cout_A31_B15, AND_A31_B15, Cout_A31_B14);

    wire AND_A0_B16;
    and and_a0_b16(AND_A0_B16, A[0], B[16]);
    wire P_A0_B16, Cout_A0_B16;
    full_adder add_a0_b16(P_A0_B16, Cout_A0_B16, P_A1_B15, AND_A0_B16, Cout_A0_B15);

    wire AND_A1_B16;
    and and_a1_b16(AND_A1_B16, A[1], B[16]);
    wire P_A1_B16, Cout_A1_B16;
    full_adder add_a1_b16(P_A1_B16, Cout_A1_B16, P_A2_B15, AND_A1_B16, Cout_A1_B15);

    wire AND_A2_B16;
    and and_a2_b16(AND_A2_B16, A[2], B[16]);
    wire P_A2_B16, Cout_A2_B16;
    full_adder add_a2_b16(P_A2_B16, Cout_A2_B16, P_A3_B15, AND_A2_B16, Cout_A2_B15);

    wire AND_A3_B16;
    and and_a3_b16(AND_A3_B16, A[3], B[16]);
    wire P_A3_B16, Cout_A3_B16;
    full_adder add_a3_b16(P_A3_B16, Cout_A3_B16, P_A4_B15, AND_A3_B16, Cout_A3_B15);

    wire AND_A4_B16;
    and and_a4_b16(AND_A4_B16, A[4], B[16]);
    wire P_A4_B16, Cout_A4_B16;
    full_adder add_a4_b16(P_A4_B16, Cout_A4_B16, P_A5_B15, AND_A4_B16, Cout_A4_B15);

    wire AND_A5_B16;
    and and_a5_b16(AND_A5_B16, A[5], B[16]);
    wire P_A5_B16, Cout_A5_B16;
    full_adder add_a5_b16(P_A5_B16, Cout_A5_B16, P_A6_B15, AND_A5_B16, Cout_A5_B15);

    wire AND_A6_B16;
    and and_a6_b16(AND_A6_B16, A[6], B[16]);
    wire P_A6_B16, Cout_A6_B16;
    full_adder add_a6_b16(P_A6_B16, Cout_A6_B16, P_A7_B15, AND_A6_B16, Cout_A6_B15);

    wire AND_A7_B16;
    and and_a7_b16(AND_A7_B16, A[7], B[16]);
    wire P_A7_B16, Cout_A7_B16;
    full_adder add_a7_b16(P_A7_B16, Cout_A7_B16, P_A8_B15, AND_A7_B16, Cout_A7_B15);

    wire AND_A8_B16;
    and and_a8_b16(AND_A8_B16, A[8], B[16]);
    wire P_A8_B16, Cout_A8_B16;
    full_adder add_a8_b16(P_A8_B16, Cout_A8_B16, P_A9_B15, AND_A8_B16, Cout_A8_B15);

    wire AND_A9_B16;
    and and_a9_b16(AND_A9_B16, A[9], B[16]);
    wire P_A9_B16, Cout_A9_B16;
    full_adder add_a9_b16(P_A9_B16, Cout_A9_B16, P_A10_B15, AND_A9_B16, Cout_A9_B15);

    wire AND_A10_B16;
    and and_a10_b16(AND_A10_B16, A[10], B[16]);
    wire P_A10_B16, Cout_A10_B16;
    full_adder add_a10_b16(P_A10_B16, Cout_A10_B16, P_A11_B15, AND_A10_B16, Cout_A10_B15);

    wire AND_A11_B16;
    and and_a11_b16(AND_A11_B16, A[11], B[16]);
    wire P_A11_B16, Cout_A11_B16;
    full_adder add_a11_b16(P_A11_B16, Cout_A11_B16, P_A12_B15, AND_A11_B16, Cout_A11_B15);

    wire AND_A12_B16;
    and and_a12_b16(AND_A12_B16, A[12], B[16]);
    wire P_A12_B16, Cout_A12_B16;
    full_adder add_a12_b16(P_A12_B16, Cout_A12_B16, P_A13_B15, AND_A12_B16, Cout_A12_B15);

    wire AND_A13_B16;
    and and_a13_b16(AND_A13_B16, A[13], B[16]);
    wire P_A13_B16, Cout_A13_B16;
    full_adder add_a13_b16(P_A13_B16, Cout_A13_B16, P_A14_B15, AND_A13_B16, Cout_A13_B15);

    wire AND_A14_B16;
    and and_a14_b16(AND_A14_B16, A[14], B[16]);
    wire P_A14_B16, Cout_A14_B16;
    full_adder add_a14_b16(P_A14_B16, Cout_A14_B16, P_A15_B15, AND_A14_B16, Cout_A14_B15);

    wire AND_A15_B16;
    and and_a15_b16(AND_A15_B16, A[15], B[16]);
    wire P_A15_B16, Cout_A15_B16;
    full_adder add_a15_b16(P_A15_B16, Cout_A15_B16, P_A16_B15, AND_A15_B16, Cout_A15_B15);

    wire AND_A16_B16;
    and and_a16_b16(AND_A16_B16, A[16], B[16]);
    wire P_A16_B16, Cout_A16_B16;
    full_adder add_a16_b16(P_A16_B16, Cout_A16_B16, P_A17_B15, AND_A16_B16, Cout_A16_B15);

    wire AND_A17_B16;
    and and_a17_b16(AND_A17_B16, A[17], B[16]);
    wire P_A17_B16, Cout_A17_B16;
    full_adder add_a17_b16(P_A17_B16, Cout_A17_B16, P_A18_B15, AND_A17_B16, Cout_A17_B15);

    wire AND_A18_B16;
    and and_a18_b16(AND_A18_B16, A[18], B[16]);
    wire P_A18_B16, Cout_A18_B16;
    full_adder add_a18_b16(P_A18_B16, Cout_A18_B16, P_A19_B15, AND_A18_B16, Cout_A18_B15);

    wire AND_A19_B16;
    and and_a19_b16(AND_A19_B16, A[19], B[16]);
    wire P_A19_B16, Cout_A19_B16;
    full_adder add_a19_b16(P_A19_B16, Cout_A19_B16, P_A20_B15, AND_A19_B16, Cout_A19_B15);

    wire AND_A20_B16;
    and and_a20_b16(AND_A20_B16, A[20], B[16]);
    wire P_A20_B16, Cout_A20_B16;
    full_adder add_a20_b16(P_A20_B16, Cout_A20_B16, P_A21_B15, AND_A20_B16, Cout_A20_B15);

    wire AND_A21_B16;
    and and_a21_b16(AND_A21_B16, A[21], B[16]);
    wire P_A21_B16, Cout_A21_B16;
    full_adder add_a21_b16(P_A21_B16, Cout_A21_B16, P_A22_B15, AND_A21_B16, Cout_A21_B15);

    wire AND_A22_B16;
    and and_a22_b16(AND_A22_B16, A[22], B[16]);
    wire P_A22_B16, Cout_A22_B16;
    full_adder add_a22_b16(P_A22_B16, Cout_A22_B16, P_A23_B15, AND_A22_B16, Cout_A22_B15);

    wire AND_A23_B16;
    and and_a23_b16(AND_A23_B16, A[23], B[16]);
    wire P_A23_B16, Cout_A23_B16;
    full_adder add_a23_b16(P_A23_B16, Cout_A23_B16, P_A24_B15, AND_A23_B16, Cout_A23_B15);

    wire AND_A24_B16;
    and and_a24_b16(AND_A24_B16, A[24], B[16]);
    wire P_A24_B16, Cout_A24_B16;
    full_adder add_a24_b16(P_A24_B16, Cout_A24_B16, P_A25_B15, AND_A24_B16, Cout_A24_B15);

    wire AND_A25_B16;
    and and_a25_b16(AND_A25_B16, A[25], B[16]);
    wire P_A25_B16, Cout_A25_B16;
    full_adder add_a25_b16(P_A25_B16, Cout_A25_B16, P_A26_B15, AND_A25_B16, Cout_A25_B15);

    wire AND_A26_B16;
    and and_a26_b16(AND_A26_B16, A[26], B[16]);
    wire P_A26_B16, Cout_A26_B16;
    full_adder add_a26_b16(P_A26_B16, Cout_A26_B16, P_A27_B15, AND_A26_B16, Cout_A26_B15);

    wire AND_A27_B16;
    and and_a27_b16(AND_A27_B16, A[27], B[16]);
    wire P_A27_B16, Cout_A27_B16;
    full_adder add_a27_b16(P_A27_B16, Cout_A27_B16, P_A28_B15, AND_A27_B16, Cout_A27_B15);

    wire AND_A28_B16;
    and and_a28_b16(AND_A28_B16, A[28], B[16]);
    wire P_A28_B16, Cout_A28_B16;
    full_adder add_a28_b16(P_A28_B16, Cout_A28_B16, P_A29_B15, AND_A28_B16, Cout_A28_B15);

    wire AND_A29_B16;
    and and_a29_b16(AND_A29_B16, A[29], B[16]);
    wire P_A29_B16, Cout_A29_B16;
    full_adder add_a29_b16(P_A29_B16, Cout_A29_B16, P_A30_B15, AND_A29_B16, Cout_A29_B15);

    wire AND_A30_B16;
    and and_a30_b16(AND_A30_B16, A[30], B[16]);
    wire P_A30_B16, Cout_A30_B16;
    full_adder add_a30_b16(P_A30_B16, Cout_A30_B16, P_A31_B15, AND_A30_B16, Cout_A30_B15);

    wire AND_A31_B16;
    nand and_a31_b16(AND_A31_B16, A[31], B[16]);
    wire P_A31_B16, Cout_A31_B16;
    half_adder add_a31_b16(P_A31_B16, Cout_A31_B16, AND_A31_B16, Cout_A31_B15);

    wire AND_A0_B17;
    and and_a0_b17(AND_A0_B17, A[0], B[17]);
    wire P_A0_B17, Cout_A0_B17;
    full_adder add_a0_b17(P_A0_B17, Cout_A0_B17, P_A1_B16, AND_A0_B17, Cout_A0_B16);

    wire AND_A1_B17;
    and and_a1_b17(AND_A1_B17, A[1], B[17]);
    wire P_A1_B17, Cout_A1_B17;
    full_adder add_a1_b17(P_A1_B17, Cout_A1_B17, P_A2_B16, AND_A1_B17, Cout_A1_B16);

    wire AND_A2_B17;
    and and_a2_b17(AND_A2_B17, A[2], B[17]);
    wire P_A2_B17, Cout_A2_B17;
    full_adder add_a2_b17(P_A2_B17, Cout_A2_B17, P_A3_B16, AND_A2_B17, Cout_A2_B16);

    wire AND_A3_B17;
    and and_a3_b17(AND_A3_B17, A[3], B[17]);
    wire P_A3_B17, Cout_A3_B17;
    full_adder add_a3_b17(P_A3_B17, Cout_A3_B17, P_A4_B16, AND_A3_B17, Cout_A3_B16);

    wire AND_A4_B17;
    and and_a4_b17(AND_A4_B17, A[4], B[17]);
    wire P_A4_B17, Cout_A4_B17;
    full_adder add_a4_b17(P_A4_B17, Cout_A4_B17, P_A5_B16, AND_A4_B17, Cout_A4_B16);

    wire AND_A5_B17;
    and and_a5_b17(AND_A5_B17, A[5], B[17]);
    wire P_A5_B17, Cout_A5_B17;
    full_adder add_a5_b17(P_A5_B17, Cout_A5_B17, P_A6_B16, AND_A5_B17, Cout_A5_B16);

    wire AND_A6_B17;
    and and_a6_b17(AND_A6_B17, A[6], B[17]);
    wire P_A6_B17, Cout_A6_B17;
    full_adder add_a6_b17(P_A6_B17, Cout_A6_B17, P_A7_B16, AND_A6_B17, Cout_A6_B16);

    wire AND_A7_B17;
    and and_a7_b17(AND_A7_B17, A[7], B[17]);
    wire P_A7_B17, Cout_A7_B17;
    full_adder add_a7_b17(P_A7_B17, Cout_A7_B17, P_A8_B16, AND_A7_B17, Cout_A7_B16);

    wire AND_A8_B17;
    and and_a8_b17(AND_A8_B17, A[8], B[17]);
    wire P_A8_B17, Cout_A8_B17;
    full_adder add_a8_b17(P_A8_B17, Cout_A8_B17, P_A9_B16, AND_A8_B17, Cout_A8_B16);

    wire AND_A9_B17;
    and and_a9_b17(AND_A9_B17, A[9], B[17]);
    wire P_A9_B17, Cout_A9_B17;
    full_adder add_a9_b17(P_A9_B17, Cout_A9_B17, P_A10_B16, AND_A9_B17, Cout_A9_B16);

    wire AND_A10_B17;
    and and_a10_b17(AND_A10_B17, A[10], B[17]);
    wire P_A10_B17, Cout_A10_B17;
    full_adder add_a10_b17(P_A10_B17, Cout_A10_B17, P_A11_B16, AND_A10_B17, Cout_A10_B16);

    wire AND_A11_B17;
    and and_a11_b17(AND_A11_B17, A[11], B[17]);
    wire P_A11_B17, Cout_A11_B17;
    full_adder add_a11_b17(P_A11_B17, Cout_A11_B17, P_A12_B16, AND_A11_B17, Cout_A11_B16);

    wire AND_A12_B17;
    and and_a12_b17(AND_A12_B17, A[12], B[17]);
    wire P_A12_B17, Cout_A12_B17;
    full_adder add_a12_b17(P_A12_B17, Cout_A12_B17, P_A13_B16, AND_A12_B17, Cout_A12_B16);

    wire AND_A13_B17;
    and and_a13_b17(AND_A13_B17, A[13], B[17]);
    wire P_A13_B17, Cout_A13_B17;
    full_adder add_a13_b17(P_A13_B17, Cout_A13_B17, P_A14_B16, AND_A13_B17, Cout_A13_B16);

    wire AND_A14_B17;
    and and_a14_b17(AND_A14_B17, A[14], B[17]);
    wire P_A14_B17, Cout_A14_B17;
    full_adder add_a14_b17(P_A14_B17, Cout_A14_B17, P_A15_B16, AND_A14_B17, Cout_A14_B16);

    wire AND_A15_B17;
    and and_a15_b17(AND_A15_B17, A[15], B[17]);
    wire P_A15_B17, Cout_A15_B17;
    full_adder add_a15_b17(P_A15_B17, Cout_A15_B17, P_A16_B16, AND_A15_B17, Cout_A15_B16);

    wire AND_A16_B17;
    and and_a16_b17(AND_A16_B17, A[16], B[17]);
    wire P_A16_B17, Cout_A16_B17;
    full_adder add_a16_b17(P_A16_B17, Cout_A16_B17, P_A17_B16, AND_A16_B17, Cout_A16_B16);

    wire AND_A17_B17;
    and and_a17_b17(AND_A17_B17, A[17], B[17]);
    wire P_A17_B17, Cout_A17_B17;
    full_adder add_a17_b17(P_A17_B17, Cout_A17_B17, P_A18_B16, AND_A17_B17, Cout_A17_B16);

    wire AND_A18_B17;
    and and_a18_b17(AND_A18_B17, A[18], B[17]);
    wire P_A18_B17, Cout_A18_B17;
    full_adder add_a18_b17(P_A18_B17, Cout_A18_B17, P_A19_B16, AND_A18_B17, Cout_A18_B16);

    wire AND_A19_B17;
    and and_a19_b17(AND_A19_B17, A[19], B[17]);
    wire P_A19_B17, Cout_A19_B17;
    full_adder add_a19_b17(P_A19_B17, Cout_A19_B17, P_A20_B16, AND_A19_B17, Cout_A19_B16);

    wire AND_A20_B17;
    and and_a20_b17(AND_A20_B17, A[20], B[17]);
    wire P_A20_B17, Cout_A20_B17;
    full_adder add_a20_b17(P_A20_B17, Cout_A20_B17, P_A21_B16, AND_A20_B17, Cout_A20_B16);

    wire AND_A21_B17;
    and and_a21_b17(AND_A21_B17, A[21], B[17]);
    wire P_A21_B17, Cout_A21_B17;
    full_adder add_a21_b17(P_A21_B17, Cout_A21_B17, P_A22_B16, AND_A21_B17, Cout_A21_B16);

    wire AND_A22_B17;
    and and_a22_b17(AND_A22_B17, A[22], B[17]);
    wire P_A22_B17, Cout_A22_B17;
    full_adder add_a22_b17(P_A22_B17, Cout_A22_B17, P_A23_B16, AND_A22_B17, Cout_A22_B16);

    wire AND_A23_B17;
    and and_a23_b17(AND_A23_B17, A[23], B[17]);
    wire P_A23_B17, Cout_A23_B17;
    full_adder add_a23_b17(P_A23_B17, Cout_A23_B17, P_A24_B16, AND_A23_B17, Cout_A23_B16);

    wire AND_A24_B17;
    and and_a24_b17(AND_A24_B17, A[24], B[17]);
    wire P_A24_B17, Cout_A24_B17;
    full_adder add_a24_b17(P_A24_B17, Cout_A24_B17, P_A25_B16, AND_A24_B17, Cout_A24_B16);

    wire AND_A25_B17;
    and and_a25_b17(AND_A25_B17, A[25], B[17]);
    wire P_A25_B17, Cout_A25_B17;
    full_adder add_a25_b17(P_A25_B17, Cout_A25_B17, P_A26_B16, AND_A25_B17, Cout_A25_B16);

    wire AND_A26_B17;
    and and_a26_b17(AND_A26_B17, A[26], B[17]);
    wire P_A26_B17, Cout_A26_B17;
    full_adder add_a26_b17(P_A26_B17, Cout_A26_B17, P_A27_B16, AND_A26_B17, Cout_A26_B16);

    wire AND_A27_B17;
    and and_a27_b17(AND_A27_B17, A[27], B[17]);
    wire P_A27_B17, Cout_A27_B17;
    full_adder add_a27_b17(P_A27_B17, Cout_A27_B17, P_A28_B16, AND_A27_B17, Cout_A27_B16);

    wire AND_A28_B17;
    and and_a28_b17(AND_A28_B17, A[28], B[17]);
    wire P_A28_B17, Cout_A28_B17;
    full_adder add_a28_b17(P_A28_B17, Cout_A28_B17, P_A29_B16, AND_A28_B17, Cout_A28_B16);

    wire AND_A29_B17;
    and and_a29_b17(AND_A29_B17, A[29], B[17]);
    wire P_A29_B17, Cout_A29_B17;
    full_adder add_a29_b17(P_A29_B17, Cout_A29_B17, P_A30_B16, AND_A29_B17, Cout_A29_B16);

    wire AND_A30_B17;
    and and_a30_b17(AND_A30_B17, A[30], B[17]);
    wire P_A30_B17, Cout_A30_B17;
    full_adder add_a30_b17(P_A30_B17, Cout_A30_B17, P_A31_B16, AND_A30_B17, Cout_A30_B16);

    wire AND_A31_B17;
    nand and_a31_b17(AND_A31_B17, A[31], B[17]);
    wire P_A31_B17, Cout_A31_B17;
    half_adder add_a31_b17(P_A31_B17, Cout_A31_B17, AND_A31_B17, Cout_A31_B16);

    wire AND_A0_B18;
    and and_a0_b18(AND_A0_B18, A[0], B[18]);
    wire P_A0_B18, Cout_A0_B18;
    full_adder add_a0_b18(P_A0_B18, Cout_A0_B18, P_A1_B17, AND_A0_B18, Cout_A0_B17);

    wire AND_A1_B18;
    and and_a1_b18(AND_A1_B18, A[1], B[18]);
    wire P_A1_B18, Cout_A1_B18;
    full_adder add_a1_b18(P_A1_B18, Cout_A1_B18, P_A2_B17, AND_A1_B18, Cout_A1_B17);

    wire AND_A2_B18;
    and and_a2_b18(AND_A2_B18, A[2], B[18]);
    wire P_A2_B18, Cout_A2_B18;
    full_adder add_a2_b18(P_A2_B18, Cout_A2_B18, P_A3_B17, AND_A2_B18, Cout_A2_B17);

    wire AND_A3_B18;
    and and_a3_b18(AND_A3_B18, A[3], B[18]);
    wire P_A3_B18, Cout_A3_B18;
    full_adder add_a3_b18(P_A3_B18, Cout_A3_B18, P_A4_B17, AND_A3_B18, Cout_A3_B17);

    wire AND_A4_B18;
    and and_a4_b18(AND_A4_B18, A[4], B[18]);
    wire P_A4_B18, Cout_A4_B18;
    full_adder add_a4_b18(P_A4_B18, Cout_A4_B18, P_A5_B17, AND_A4_B18, Cout_A4_B17);

    wire AND_A5_B18;
    and and_a5_b18(AND_A5_B18, A[5], B[18]);
    wire P_A5_B18, Cout_A5_B18;
    full_adder add_a5_b18(P_A5_B18, Cout_A5_B18, P_A6_B17, AND_A5_B18, Cout_A5_B17);

    wire AND_A6_B18;
    and and_a6_b18(AND_A6_B18, A[6], B[18]);
    wire P_A6_B18, Cout_A6_B18;
    full_adder add_a6_b18(P_A6_B18, Cout_A6_B18, P_A7_B17, AND_A6_B18, Cout_A6_B17);

    wire AND_A7_B18;
    and and_a7_b18(AND_A7_B18, A[7], B[18]);
    wire P_A7_B18, Cout_A7_B18;
    full_adder add_a7_b18(P_A7_B18, Cout_A7_B18, P_A8_B17, AND_A7_B18, Cout_A7_B17);

    wire AND_A8_B18;
    and and_a8_b18(AND_A8_B18, A[8], B[18]);
    wire P_A8_B18, Cout_A8_B18;
    full_adder add_a8_b18(P_A8_B18, Cout_A8_B18, P_A9_B17, AND_A8_B18, Cout_A8_B17);

    wire AND_A9_B18;
    and and_a9_b18(AND_A9_B18, A[9], B[18]);
    wire P_A9_B18, Cout_A9_B18;
    full_adder add_a9_b18(P_A9_B18, Cout_A9_B18, P_A10_B17, AND_A9_B18, Cout_A9_B17);

    wire AND_A10_B18;
    and and_a10_b18(AND_A10_B18, A[10], B[18]);
    wire P_A10_B18, Cout_A10_B18;
    full_adder add_a10_b18(P_A10_B18, Cout_A10_B18, P_A11_B17, AND_A10_B18, Cout_A10_B17);

    wire AND_A11_B18;
    and and_a11_b18(AND_A11_B18, A[11], B[18]);
    wire P_A11_B18, Cout_A11_B18;
    full_adder add_a11_b18(P_A11_B18, Cout_A11_B18, P_A12_B17, AND_A11_B18, Cout_A11_B17);

    wire AND_A12_B18;
    and and_a12_b18(AND_A12_B18, A[12], B[18]);
    wire P_A12_B18, Cout_A12_B18;
    full_adder add_a12_b18(P_A12_B18, Cout_A12_B18, P_A13_B17, AND_A12_B18, Cout_A12_B17);

    wire AND_A13_B18;
    and and_a13_b18(AND_A13_B18, A[13], B[18]);
    wire P_A13_B18, Cout_A13_B18;
    full_adder add_a13_b18(P_A13_B18, Cout_A13_B18, P_A14_B17, AND_A13_B18, Cout_A13_B17);

    wire AND_A14_B18;
    and and_a14_b18(AND_A14_B18, A[14], B[18]);
    wire P_A14_B18, Cout_A14_B18;
    full_adder add_a14_b18(P_A14_B18, Cout_A14_B18, P_A15_B17, AND_A14_B18, Cout_A14_B17);

    wire AND_A15_B18;
    and and_a15_b18(AND_A15_B18, A[15], B[18]);
    wire P_A15_B18, Cout_A15_B18;
    full_adder add_a15_b18(P_A15_B18, Cout_A15_B18, P_A16_B17, AND_A15_B18, Cout_A15_B17);

    wire AND_A16_B18;
    and and_a16_b18(AND_A16_B18, A[16], B[18]);
    wire P_A16_B18, Cout_A16_B18;
    full_adder add_a16_b18(P_A16_B18, Cout_A16_B18, P_A17_B17, AND_A16_B18, Cout_A16_B17);

    wire AND_A17_B18;
    and and_a17_b18(AND_A17_B18, A[17], B[18]);
    wire P_A17_B18, Cout_A17_B18;
    full_adder add_a17_b18(P_A17_B18, Cout_A17_B18, P_A18_B17, AND_A17_B18, Cout_A17_B17);

    wire AND_A18_B18;
    and and_a18_b18(AND_A18_B18, A[18], B[18]);
    wire P_A18_B18, Cout_A18_B18;
    full_adder add_a18_b18(P_A18_B18, Cout_A18_B18, P_A19_B17, AND_A18_B18, Cout_A18_B17);

    wire AND_A19_B18;
    and and_a19_b18(AND_A19_B18, A[19], B[18]);
    wire P_A19_B18, Cout_A19_B18;
    full_adder add_a19_b18(P_A19_B18, Cout_A19_B18, P_A20_B17, AND_A19_B18, Cout_A19_B17);

    wire AND_A20_B18;
    and and_a20_b18(AND_A20_B18, A[20], B[18]);
    wire P_A20_B18, Cout_A20_B18;
    full_adder add_a20_b18(P_A20_B18, Cout_A20_B18, P_A21_B17, AND_A20_B18, Cout_A20_B17);

    wire AND_A21_B18;
    and and_a21_b18(AND_A21_B18, A[21], B[18]);
    wire P_A21_B18, Cout_A21_B18;
    full_adder add_a21_b18(P_A21_B18, Cout_A21_B18, P_A22_B17, AND_A21_B18, Cout_A21_B17);

    wire AND_A22_B18;
    and and_a22_b18(AND_A22_B18, A[22], B[18]);
    wire P_A22_B18, Cout_A22_B18;
    full_adder add_a22_b18(P_A22_B18, Cout_A22_B18, P_A23_B17, AND_A22_B18, Cout_A22_B17);

    wire AND_A23_B18;
    and and_a23_b18(AND_A23_B18, A[23], B[18]);
    wire P_A23_B18, Cout_A23_B18;
    full_adder add_a23_b18(P_A23_B18, Cout_A23_B18, P_A24_B17, AND_A23_B18, Cout_A23_B17);

    wire AND_A24_B18;
    and and_a24_b18(AND_A24_B18, A[24], B[18]);
    wire P_A24_B18, Cout_A24_B18;
    full_adder add_a24_b18(P_A24_B18, Cout_A24_B18, P_A25_B17, AND_A24_B18, Cout_A24_B17);

    wire AND_A25_B18;
    and and_a25_b18(AND_A25_B18, A[25], B[18]);
    wire P_A25_B18, Cout_A25_B18;
    full_adder add_a25_b18(P_A25_B18, Cout_A25_B18, P_A26_B17, AND_A25_B18, Cout_A25_B17);

    wire AND_A26_B18;
    and and_a26_b18(AND_A26_B18, A[26], B[18]);
    wire P_A26_B18, Cout_A26_B18;
    full_adder add_a26_b18(P_A26_B18, Cout_A26_B18, P_A27_B17, AND_A26_B18, Cout_A26_B17);

    wire AND_A27_B18;
    and and_a27_b18(AND_A27_B18, A[27], B[18]);
    wire P_A27_B18, Cout_A27_B18;
    full_adder add_a27_b18(P_A27_B18, Cout_A27_B18, P_A28_B17, AND_A27_B18, Cout_A27_B17);

    wire AND_A28_B18;
    and and_a28_b18(AND_A28_B18, A[28], B[18]);
    wire P_A28_B18, Cout_A28_B18;
    full_adder add_a28_b18(P_A28_B18, Cout_A28_B18, P_A29_B17, AND_A28_B18, Cout_A28_B17);

    wire AND_A29_B18;
    and and_a29_b18(AND_A29_B18, A[29], B[18]);
    wire P_A29_B18, Cout_A29_B18;
    full_adder add_a29_b18(P_A29_B18, Cout_A29_B18, P_A30_B17, AND_A29_B18, Cout_A29_B17);

    wire AND_A30_B18;
    and and_a30_b18(AND_A30_B18, A[30], B[18]);
    wire P_A30_B18, Cout_A30_B18;
    full_adder add_a30_b18(P_A30_B18, Cout_A30_B18, P_A31_B17, AND_A30_B18, Cout_A30_B17);

    wire AND_A31_B18;
    nand and_a31_b18(AND_A31_B18, A[31], B[18]);
    wire P_A31_B18, Cout_A31_B18;
    half_adder add_a31_b18(P_A31_B18, Cout_A31_B18, AND_A31_B18, Cout_A31_B17);

    wire AND_A0_B19;
    and and_a0_b19(AND_A0_B19, A[0], B[19]);
    wire P_A0_B19, Cout_A0_B19;
    full_adder add_a0_b19(P_A0_B19, Cout_A0_B19, P_A1_B18, AND_A0_B19, Cout_A0_B18);

    wire AND_A1_B19;
    and and_a1_b19(AND_A1_B19, A[1], B[19]);
    wire P_A1_B19, Cout_A1_B19;
    full_adder add_a1_b19(P_A1_B19, Cout_A1_B19, P_A2_B18, AND_A1_B19, Cout_A1_B18);

    wire AND_A2_B19;
    and and_a2_b19(AND_A2_B19, A[2], B[19]);
    wire P_A2_B19, Cout_A2_B19;
    full_adder add_a2_b19(P_A2_B19, Cout_A2_B19, P_A3_B18, AND_A2_B19, Cout_A2_B18);

    wire AND_A3_B19;
    and and_a3_b19(AND_A3_B19, A[3], B[19]);
    wire P_A3_B19, Cout_A3_B19;
    full_adder add_a3_b19(P_A3_B19, Cout_A3_B19, P_A4_B18, AND_A3_B19, Cout_A3_B18);

    wire AND_A4_B19;
    and and_a4_b19(AND_A4_B19, A[4], B[19]);
    wire P_A4_B19, Cout_A4_B19;
    full_adder add_a4_b19(P_A4_B19, Cout_A4_B19, P_A5_B18, AND_A4_B19, Cout_A4_B18);

    wire AND_A5_B19;
    and and_a5_b19(AND_A5_B19, A[5], B[19]);
    wire P_A5_B19, Cout_A5_B19;
    full_adder add_a5_b19(P_A5_B19, Cout_A5_B19, P_A6_B18, AND_A5_B19, Cout_A5_B18);

    wire AND_A6_B19;
    and and_a6_b19(AND_A6_B19, A[6], B[19]);
    wire P_A6_B19, Cout_A6_B19;
    full_adder add_a6_b19(P_A6_B19, Cout_A6_B19, P_A7_B18, AND_A6_B19, Cout_A6_B18);

    wire AND_A7_B19;
    and and_a7_b19(AND_A7_B19, A[7], B[19]);
    wire P_A7_B19, Cout_A7_B19;
    full_adder add_a7_b19(P_A7_B19, Cout_A7_B19, P_A8_B18, AND_A7_B19, Cout_A7_B18);

    wire AND_A8_B19;
    and and_a8_b19(AND_A8_B19, A[8], B[19]);
    wire P_A8_B19, Cout_A8_B19;
    full_adder add_a8_b19(P_A8_B19, Cout_A8_B19, P_A9_B18, AND_A8_B19, Cout_A8_B18);

    wire AND_A9_B19;
    and and_a9_b19(AND_A9_B19, A[9], B[19]);
    wire P_A9_B19, Cout_A9_B19;
    full_adder add_a9_b19(P_A9_B19, Cout_A9_B19, P_A10_B18, AND_A9_B19, Cout_A9_B18);

    wire AND_A10_B19;
    and and_a10_b19(AND_A10_B19, A[10], B[19]);
    wire P_A10_B19, Cout_A10_B19;
    full_adder add_a10_b19(P_A10_B19, Cout_A10_B19, P_A11_B18, AND_A10_B19, Cout_A10_B18);

    wire AND_A11_B19;
    and and_a11_b19(AND_A11_B19, A[11], B[19]);
    wire P_A11_B19, Cout_A11_B19;
    full_adder add_a11_b19(P_A11_B19, Cout_A11_B19, P_A12_B18, AND_A11_B19, Cout_A11_B18);

    wire AND_A12_B19;
    and and_a12_b19(AND_A12_B19, A[12], B[19]);
    wire P_A12_B19, Cout_A12_B19;
    full_adder add_a12_b19(P_A12_B19, Cout_A12_B19, P_A13_B18, AND_A12_B19, Cout_A12_B18);

    wire AND_A13_B19;
    and and_a13_b19(AND_A13_B19, A[13], B[19]);
    wire P_A13_B19, Cout_A13_B19;
    full_adder add_a13_b19(P_A13_B19, Cout_A13_B19, P_A14_B18, AND_A13_B19, Cout_A13_B18);

    wire AND_A14_B19;
    and and_a14_b19(AND_A14_B19, A[14], B[19]);
    wire P_A14_B19, Cout_A14_B19;
    full_adder add_a14_b19(P_A14_B19, Cout_A14_B19, P_A15_B18, AND_A14_B19, Cout_A14_B18);

    wire AND_A15_B19;
    and and_a15_b19(AND_A15_B19, A[15], B[19]);
    wire P_A15_B19, Cout_A15_B19;
    full_adder add_a15_b19(P_A15_B19, Cout_A15_B19, P_A16_B18, AND_A15_B19, Cout_A15_B18);

    wire AND_A16_B19;
    and and_a16_b19(AND_A16_B19, A[16], B[19]);
    wire P_A16_B19, Cout_A16_B19;
    full_adder add_a16_b19(P_A16_B19, Cout_A16_B19, P_A17_B18, AND_A16_B19, Cout_A16_B18);

    wire AND_A17_B19;
    and and_a17_b19(AND_A17_B19, A[17], B[19]);
    wire P_A17_B19, Cout_A17_B19;
    full_adder add_a17_b19(P_A17_B19, Cout_A17_B19, P_A18_B18, AND_A17_B19, Cout_A17_B18);

    wire AND_A18_B19;
    and and_a18_b19(AND_A18_B19, A[18], B[19]);
    wire P_A18_B19, Cout_A18_B19;
    full_adder add_a18_b19(P_A18_B19, Cout_A18_B19, P_A19_B18, AND_A18_B19, Cout_A18_B18);

    wire AND_A19_B19;
    and and_a19_b19(AND_A19_B19, A[19], B[19]);
    wire P_A19_B19, Cout_A19_B19;
    full_adder add_a19_b19(P_A19_B19, Cout_A19_B19, P_A20_B18, AND_A19_B19, Cout_A19_B18);

    wire AND_A20_B19;
    and and_a20_b19(AND_A20_B19, A[20], B[19]);
    wire P_A20_B19, Cout_A20_B19;
    full_adder add_a20_b19(P_A20_B19, Cout_A20_B19, P_A21_B18, AND_A20_B19, Cout_A20_B18);

    wire AND_A21_B19;
    and and_a21_b19(AND_A21_B19, A[21], B[19]);
    wire P_A21_B19, Cout_A21_B19;
    full_adder add_a21_b19(P_A21_B19, Cout_A21_B19, P_A22_B18, AND_A21_B19, Cout_A21_B18);

    wire AND_A22_B19;
    and and_a22_b19(AND_A22_B19, A[22], B[19]);
    wire P_A22_B19, Cout_A22_B19;
    full_adder add_a22_b19(P_A22_B19, Cout_A22_B19, P_A23_B18, AND_A22_B19, Cout_A22_B18);

    wire AND_A23_B19;
    and and_a23_b19(AND_A23_B19, A[23], B[19]);
    wire P_A23_B19, Cout_A23_B19;
    full_adder add_a23_b19(P_A23_B19, Cout_A23_B19, P_A24_B18, AND_A23_B19, Cout_A23_B18);

    wire AND_A24_B19;
    and and_a24_b19(AND_A24_B19, A[24], B[19]);
    wire P_A24_B19, Cout_A24_B19;
    full_adder add_a24_b19(P_A24_B19, Cout_A24_B19, P_A25_B18, AND_A24_B19, Cout_A24_B18);

    wire AND_A25_B19;
    and and_a25_b19(AND_A25_B19, A[25], B[19]);
    wire P_A25_B19, Cout_A25_B19;
    full_adder add_a25_b19(P_A25_B19, Cout_A25_B19, P_A26_B18, AND_A25_B19, Cout_A25_B18);

    wire AND_A26_B19;
    and and_a26_b19(AND_A26_B19, A[26], B[19]);
    wire P_A26_B19, Cout_A26_B19;
    full_adder add_a26_b19(P_A26_B19, Cout_A26_B19, P_A27_B18, AND_A26_B19, Cout_A26_B18);

    wire AND_A27_B19;
    and and_a27_b19(AND_A27_B19, A[27], B[19]);
    wire P_A27_B19, Cout_A27_B19;
    full_adder add_a27_b19(P_A27_B19, Cout_A27_B19, P_A28_B18, AND_A27_B19, Cout_A27_B18);

    wire AND_A28_B19;
    and and_a28_b19(AND_A28_B19, A[28], B[19]);
    wire P_A28_B19, Cout_A28_B19;
    full_adder add_a28_b19(P_A28_B19, Cout_A28_B19, P_A29_B18, AND_A28_B19, Cout_A28_B18);

    wire AND_A29_B19;
    and and_a29_b19(AND_A29_B19, A[29], B[19]);
    wire P_A29_B19, Cout_A29_B19;
    full_adder add_a29_b19(P_A29_B19, Cout_A29_B19, P_A30_B18, AND_A29_B19, Cout_A29_B18);

    wire AND_A30_B19;
    and and_a30_b19(AND_A30_B19, A[30], B[19]);
    wire P_A30_B19, Cout_A30_B19;
    full_adder add_a30_b19(P_A30_B19, Cout_A30_B19, P_A31_B18, AND_A30_B19, Cout_A30_B18);

    wire AND_A31_B19;
    nand and_a31_b19(AND_A31_B19, A[31], B[19]);
    wire P_A31_B19, Cout_A31_B19;
    half_adder add_a31_b19(P_A31_B19, Cout_A31_B19, AND_A31_B19, Cout_A31_B18);

    wire AND_A0_B20;
    and and_a0_b20(AND_A0_B20, A[0], B[20]);
    wire P_A0_B20, Cout_A0_B20;
    full_adder add_a0_b20(P_A0_B20, Cout_A0_B20, P_A1_B19, AND_A0_B20, Cout_A0_B19);

    wire AND_A1_B20;
    and and_a1_b20(AND_A1_B20, A[1], B[20]);
    wire P_A1_B20, Cout_A1_B20;
    full_adder add_a1_b20(P_A1_B20, Cout_A1_B20, P_A2_B19, AND_A1_B20, Cout_A1_B19);

    wire AND_A2_B20;
    and and_a2_b20(AND_A2_B20, A[2], B[20]);
    wire P_A2_B20, Cout_A2_B20;
    full_adder add_a2_b20(P_A2_B20, Cout_A2_B20, P_A3_B19, AND_A2_B20, Cout_A2_B19);

    wire AND_A3_B20;
    and and_a3_b20(AND_A3_B20, A[3], B[20]);
    wire P_A3_B20, Cout_A3_B20;
    full_adder add_a3_b20(P_A3_B20, Cout_A3_B20, P_A4_B19, AND_A3_B20, Cout_A3_B19);

    wire AND_A4_B20;
    and and_a4_b20(AND_A4_B20, A[4], B[20]);
    wire P_A4_B20, Cout_A4_B20;
    full_adder add_a4_b20(P_A4_B20, Cout_A4_B20, P_A5_B19, AND_A4_B20, Cout_A4_B19);

    wire AND_A5_B20;
    and and_a5_b20(AND_A5_B20, A[5], B[20]);
    wire P_A5_B20, Cout_A5_B20;
    full_adder add_a5_b20(P_A5_B20, Cout_A5_B20, P_A6_B19, AND_A5_B20, Cout_A5_B19);

    wire AND_A6_B20;
    and and_a6_b20(AND_A6_B20, A[6], B[20]);
    wire P_A6_B20, Cout_A6_B20;
    full_adder add_a6_b20(P_A6_B20, Cout_A6_B20, P_A7_B19, AND_A6_B20, Cout_A6_B19);

    wire AND_A7_B20;
    and and_a7_b20(AND_A7_B20, A[7], B[20]);
    wire P_A7_B20, Cout_A7_B20;
    full_adder add_a7_b20(P_A7_B20, Cout_A7_B20, P_A8_B19, AND_A7_B20, Cout_A7_B19);

    wire AND_A8_B20;
    and and_a8_b20(AND_A8_B20, A[8], B[20]);
    wire P_A8_B20, Cout_A8_B20;
    full_adder add_a8_b20(P_A8_B20, Cout_A8_B20, P_A9_B19, AND_A8_B20, Cout_A8_B19);

    wire AND_A9_B20;
    and and_a9_b20(AND_A9_B20, A[9], B[20]);
    wire P_A9_B20, Cout_A9_B20;
    full_adder add_a9_b20(P_A9_B20, Cout_A9_B20, P_A10_B19, AND_A9_B20, Cout_A9_B19);

    wire AND_A10_B20;
    and and_a10_b20(AND_A10_B20, A[10], B[20]);
    wire P_A10_B20, Cout_A10_B20;
    full_adder add_a10_b20(P_A10_B20, Cout_A10_B20, P_A11_B19, AND_A10_B20, Cout_A10_B19);

    wire AND_A11_B20;
    and and_a11_b20(AND_A11_B20, A[11], B[20]);
    wire P_A11_B20, Cout_A11_B20;
    full_adder add_a11_b20(P_A11_B20, Cout_A11_B20, P_A12_B19, AND_A11_B20, Cout_A11_B19);

    wire AND_A12_B20;
    and and_a12_b20(AND_A12_B20, A[12], B[20]);
    wire P_A12_B20, Cout_A12_B20;
    full_adder add_a12_b20(P_A12_B20, Cout_A12_B20, P_A13_B19, AND_A12_B20, Cout_A12_B19);

    wire AND_A13_B20;
    and and_a13_b20(AND_A13_B20, A[13], B[20]);
    wire P_A13_B20, Cout_A13_B20;
    full_adder add_a13_b20(P_A13_B20, Cout_A13_B20, P_A14_B19, AND_A13_B20, Cout_A13_B19);

    wire AND_A14_B20;
    and and_a14_b20(AND_A14_B20, A[14], B[20]);
    wire P_A14_B20, Cout_A14_B20;
    full_adder add_a14_b20(P_A14_B20, Cout_A14_B20, P_A15_B19, AND_A14_B20, Cout_A14_B19);

    wire AND_A15_B20;
    and and_a15_b20(AND_A15_B20, A[15], B[20]);
    wire P_A15_B20, Cout_A15_B20;
    full_adder add_a15_b20(P_A15_B20, Cout_A15_B20, P_A16_B19, AND_A15_B20, Cout_A15_B19);

    wire AND_A16_B20;
    and and_a16_b20(AND_A16_B20, A[16], B[20]);
    wire P_A16_B20, Cout_A16_B20;
    full_adder add_a16_b20(P_A16_B20, Cout_A16_B20, P_A17_B19, AND_A16_B20, Cout_A16_B19);

    wire AND_A17_B20;
    and and_a17_b20(AND_A17_B20, A[17], B[20]);
    wire P_A17_B20, Cout_A17_B20;
    full_adder add_a17_b20(P_A17_B20, Cout_A17_B20, P_A18_B19, AND_A17_B20, Cout_A17_B19);

    wire AND_A18_B20;
    and and_a18_b20(AND_A18_B20, A[18], B[20]);
    wire P_A18_B20, Cout_A18_B20;
    full_adder add_a18_b20(P_A18_B20, Cout_A18_B20, P_A19_B19, AND_A18_B20, Cout_A18_B19);

    wire AND_A19_B20;
    and and_a19_b20(AND_A19_B20, A[19], B[20]);
    wire P_A19_B20, Cout_A19_B20;
    full_adder add_a19_b20(P_A19_B20, Cout_A19_B20, P_A20_B19, AND_A19_B20, Cout_A19_B19);

    wire AND_A20_B20;
    and and_a20_b20(AND_A20_B20, A[20], B[20]);
    wire P_A20_B20, Cout_A20_B20;
    full_adder add_a20_b20(P_A20_B20, Cout_A20_B20, P_A21_B19, AND_A20_B20, Cout_A20_B19);

    wire AND_A21_B20;
    and and_a21_b20(AND_A21_B20, A[21], B[20]);
    wire P_A21_B20, Cout_A21_B20;
    full_adder add_a21_b20(P_A21_B20, Cout_A21_B20, P_A22_B19, AND_A21_B20, Cout_A21_B19);

    wire AND_A22_B20;
    and and_a22_b20(AND_A22_B20, A[22], B[20]);
    wire P_A22_B20, Cout_A22_B20;
    full_adder add_a22_b20(P_A22_B20, Cout_A22_B20, P_A23_B19, AND_A22_B20, Cout_A22_B19);

    wire AND_A23_B20;
    and and_a23_b20(AND_A23_B20, A[23], B[20]);
    wire P_A23_B20, Cout_A23_B20;
    full_adder add_a23_b20(P_A23_B20, Cout_A23_B20, P_A24_B19, AND_A23_B20, Cout_A23_B19);

    wire AND_A24_B20;
    and and_a24_b20(AND_A24_B20, A[24], B[20]);
    wire P_A24_B20, Cout_A24_B20;
    full_adder add_a24_b20(P_A24_B20, Cout_A24_B20, P_A25_B19, AND_A24_B20, Cout_A24_B19);

    wire AND_A25_B20;
    and and_a25_b20(AND_A25_B20, A[25], B[20]);
    wire P_A25_B20, Cout_A25_B20;
    full_adder add_a25_b20(P_A25_B20, Cout_A25_B20, P_A26_B19, AND_A25_B20, Cout_A25_B19);

    wire AND_A26_B20;
    and and_a26_b20(AND_A26_B20, A[26], B[20]);
    wire P_A26_B20, Cout_A26_B20;
    full_adder add_a26_b20(P_A26_B20, Cout_A26_B20, P_A27_B19, AND_A26_B20, Cout_A26_B19);

    wire AND_A27_B20;
    and and_a27_b20(AND_A27_B20, A[27], B[20]);
    wire P_A27_B20, Cout_A27_B20;
    full_adder add_a27_b20(P_A27_B20, Cout_A27_B20, P_A28_B19, AND_A27_B20, Cout_A27_B19);

    wire AND_A28_B20;
    and and_a28_b20(AND_A28_B20, A[28], B[20]);
    wire P_A28_B20, Cout_A28_B20;
    full_adder add_a28_b20(P_A28_B20, Cout_A28_B20, P_A29_B19, AND_A28_B20, Cout_A28_B19);

    wire AND_A29_B20;
    and and_a29_b20(AND_A29_B20, A[29], B[20]);
    wire P_A29_B20, Cout_A29_B20;
    full_adder add_a29_b20(P_A29_B20, Cout_A29_B20, P_A30_B19, AND_A29_B20, Cout_A29_B19);

    wire AND_A30_B20;
    and and_a30_b20(AND_A30_B20, A[30], B[20]);
    wire P_A30_B20, Cout_A30_B20;
    full_adder add_a30_b20(P_A30_B20, Cout_A30_B20, P_A31_B19, AND_A30_B20, Cout_A30_B19);

    wire AND_A31_B20;
    nand and_a31_b20(AND_A31_B20, A[31], B[20]);
    wire P_A31_B20, Cout_A31_B20;
    half_adder add_a31_b20(P_A31_B20, Cout_A31_B20, AND_A31_B20, Cout_A31_B19);

    wire AND_A0_B21;
    and and_a0_b21(AND_A0_B21, A[0], B[21]);
    wire P_A0_B21, Cout_A0_B21;
    full_adder add_a0_b21(P_A0_B21, Cout_A0_B21, P_A1_B20, AND_A0_B21, Cout_A0_B20);

    wire AND_A1_B21;
    and and_a1_b21(AND_A1_B21, A[1], B[21]);
    wire P_A1_B21, Cout_A1_B21;
    full_adder add_a1_b21(P_A1_B21, Cout_A1_B21, P_A2_B20, AND_A1_B21, Cout_A1_B20);

    wire AND_A2_B21;
    and and_a2_b21(AND_A2_B21, A[2], B[21]);
    wire P_A2_B21, Cout_A2_B21;
    full_adder add_a2_b21(P_A2_B21, Cout_A2_B21, P_A3_B20, AND_A2_B21, Cout_A2_B20);

    wire AND_A3_B21;
    and and_a3_b21(AND_A3_B21, A[3], B[21]);
    wire P_A3_B21, Cout_A3_B21;
    full_adder add_a3_b21(P_A3_B21, Cout_A3_B21, P_A4_B20, AND_A3_B21, Cout_A3_B20);

    wire AND_A4_B21;
    and and_a4_b21(AND_A4_B21, A[4], B[21]);
    wire P_A4_B21, Cout_A4_B21;
    full_adder add_a4_b21(P_A4_B21, Cout_A4_B21, P_A5_B20, AND_A4_B21, Cout_A4_B20);

    wire AND_A5_B21;
    and and_a5_b21(AND_A5_B21, A[5], B[21]);
    wire P_A5_B21, Cout_A5_B21;
    full_adder add_a5_b21(P_A5_B21, Cout_A5_B21, P_A6_B20, AND_A5_B21, Cout_A5_B20);

    wire AND_A6_B21;
    and and_a6_b21(AND_A6_B21, A[6], B[21]);
    wire P_A6_B21, Cout_A6_B21;
    full_adder add_a6_b21(P_A6_B21, Cout_A6_B21, P_A7_B20, AND_A6_B21, Cout_A6_B20);

    wire AND_A7_B21;
    and and_a7_b21(AND_A7_B21, A[7], B[21]);
    wire P_A7_B21, Cout_A7_B21;
    full_adder add_a7_b21(P_A7_B21, Cout_A7_B21, P_A8_B20, AND_A7_B21, Cout_A7_B20);

    wire AND_A8_B21;
    and and_a8_b21(AND_A8_B21, A[8], B[21]);
    wire P_A8_B21, Cout_A8_B21;
    full_adder add_a8_b21(P_A8_B21, Cout_A8_B21, P_A9_B20, AND_A8_B21, Cout_A8_B20);

    wire AND_A9_B21;
    and and_a9_b21(AND_A9_B21, A[9], B[21]);
    wire P_A9_B21, Cout_A9_B21;
    full_adder add_a9_b21(P_A9_B21, Cout_A9_B21, P_A10_B20, AND_A9_B21, Cout_A9_B20);

    wire AND_A10_B21;
    and and_a10_b21(AND_A10_B21, A[10], B[21]);
    wire P_A10_B21, Cout_A10_B21;
    full_adder add_a10_b21(P_A10_B21, Cout_A10_B21, P_A11_B20, AND_A10_B21, Cout_A10_B20);

    wire AND_A11_B21;
    and and_a11_b21(AND_A11_B21, A[11], B[21]);
    wire P_A11_B21, Cout_A11_B21;
    full_adder add_a11_b21(P_A11_B21, Cout_A11_B21, P_A12_B20, AND_A11_B21, Cout_A11_B20);

    wire AND_A12_B21;
    and and_a12_b21(AND_A12_B21, A[12], B[21]);
    wire P_A12_B21, Cout_A12_B21;
    full_adder add_a12_b21(P_A12_B21, Cout_A12_B21, P_A13_B20, AND_A12_B21, Cout_A12_B20);

    wire AND_A13_B21;
    and and_a13_b21(AND_A13_B21, A[13], B[21]);
    wire P_A13_B21, Cout_A13_B21;
    full_adder add_a13_b21(P_A13_B21, Cout_A13_B21, P_A14_B20, AND_A13_B21, Cout_A13_B20);

    wire AND_A14_B21;
    and and_a14_b21(AND_A14_B21, A[14], B[21]);
    wire P_A14_B21, Cout_A14_B21;
    full_adder add_a14_b21(P_A14_B21, Cout_A14_B21, P_A15_B20, AND_A14_B21, Cout_A14_B20);

    wire AND_A15_B21;
    and and_a15_b21(AND_A15_B21, A[15], B[21]);
    wire P_A15_B21, Cout_A15_B21;
    full_adder add_a15_b21(P_A15_B21, Cout_A15_B21, P_A16_B20, AND_A15_B21, Cout_A15_B20);

    wire AND_A16_B21;
    and and_a16_b21(AND_A16_B21, A[16], B[21]);
    wire P_A16_B21, Cout_A16_B21;
    full_adder add_a16_b21(P_A16_B21, Cout_A16_B21, P_A17_B20, AND_A16_B21, Cout_A16_B20);

    wire AND_A17_B21;
    and and_a17_b21(AND_A17_B21, A[17], B[21]);
    wire P_A17_B21, Cout_A17_B21;
    full_adder add_a17_b21(P_A17_B21, Cout_A17_B21, P_A18_B20, AND_A17_B21, Cout_A17_B20);

    wire AND_A18_B21;
    and and_a18_b21(AND_A18_B21, A[18], B[21]);
    wire P_A18_B21, Cout_A18_B21;
    full_adder add_a18_b21(P_A18_B21, Cout_A18_B21, P_A19_B20, AND_A18_B21, Cout_A18_B20);

    wire AND_A19_B21;
    and and_a19_b21(AND_A19_B21, A[19], B[21]);
    wire P_A19_B21, Cout_A19_B21;
    full_adder add_a19_b21(P_A19_B21, Cout_A19_B21, P_A20_B20, AND_A19_B21, Cout_A19_B20);

    wire AND_A20_B21;
    and and_a20_b21(AND_A20_B21, A[20], B[21]);
    wire P_A20_B21, Cout_A20_B21;
    full_adder add_a20_b21(P_A20_B21, Cout_A20_B21, P_A21_B20, AND_A20_B21, Cout_A20_B20);

    wire AND_A21_B21;
    and and_a21_b21(AND_A21_B21, A[21], B[21]);
    wire P_A21_B21, Cout_A21_B21;
    full_adder add_a21_b21(P_A21_B21, Cout_A21_B21, P_A22_B20, AND_A21_B21, Cout_A21_B20);

    wire AND_A22_B21;
    and and_a22_b21(AND_A22_B21, A[22], B[21]);
    wire P_A22_B21, Cout_A22_B21;
    full_adder add_a22_b21(P_A22_B21, Cout_A22_B21, P_A23_B20, AND_A22_B21, Cout_A22_B20);

    wire AND_A23_B21;
    and and_a23_b21(AND_A23_B21, A[23], B[21]);
    wire P_A23_B21, Cout_A23_B21;
    full_adder add_a23_b21(P_A23_B21, Cout_A23_B21, P_A24_B20, AND_A23_B21, Cout_A23_B20);

    wire AND_A24_B21;
    and and_a24_b21(AND_A24_B21, A[24], B[21]);
    wire P_A24_B21, Cout_A24_B21;
    full_adder add_a24_b21(P_A24_B21, Cout_A24_B21, P_A25_B20, AND_A24_B21, Cout_A24_B20);

    wire AND_A25_B21;
    and and_a25_b21(AND_A25_B21, A[25], B[21]);
    wire P_A25_B21, Cout_A25_B21;
    full_adder add_a25_b21(P_A25_B21, Cout_A25_B21, P_A26_B20, AND_A25_B21, Cout_A25_B20);

    wire AND_A26_B21;
    and and_a26_b21(AND_A26_B21, A[26], B[21]);
    wire P_A26_B21, Cout_A26_B21;
    full_adder add_a26_b21(P_A26_B21, Cout_A26_B21, P_A27_B20, AND_A26_B21, Cout_A26_B20);

    wire AND_A27_B21;
    and and_a27_b21(AND_A27_B21, A[27], B[21]);
    wire P_A27_B21, Cout_A27_B21;
    full_adder add_a27_b21(P_A27_B21, Cout_A27_B21, P_A28_B20, AND_A27_B21, Cout_A27_B20);

    wire AND_A28_B21;
    and and_a28_b21(AND_A28_B21, A[28], B[21]);
    wire P_A28_B21, Cout_A28_B21;
    full_adder add_a28_b21(P_A28_B21, Cout_A28_B21, P_A29_B20, AND_A28_B21, Cout_A28_B20);

    wire AND_A29_B21;
    and and_a29_b21(AND_A29_B21, A[29], B[21]);
    wire P_A29_B21, Cout_A29_B21;
    full_adder add_a29_b21(P_A29_B21, Cout_A29_B21, P_A30_B20, AND_A29_B21, Cout_A29_B20);

    wire AND_A30_B21;
    and and_a30_b21(AND_A30_B21, A[30], B[21]);
    wire P_A30_B21, Cout_A30_B21;
    full_adder add_a30_b21(P_A30_B21, Cout_A30_B21, P_A31_B20, AND_A30_B21, Cout_A30_B20);

    wire AND_A31_B21;
    nand and_a31_b21(AND_A31_B21, A[31], B[21]);
    wire P_A31_B21, Cout_A31_B21;
    half_adder add_a31_b21(P_A31_B21, Cout_A31_B21, AND_A31_B21, Cout_A31_B20);

    wire AND_A0_B22;
    and and_a0_b22(AND_A0_B22, A[0], B[22]);
    wire P_A0_B22, Cout_A0_B22;
    full_adder add_a0_b22(P_A0_B22, Cout_A0_B22, P_A1_B21, AND_A0_B22, Cout_A0_B21);

    wire AND_A1_B22;
    and and_a1_b22(AND_A1_B22, A[1], B[22]);
    wire P_A1_B22, Cout_A1_B22;
    full_adder add_a1_b22(P_A1_B22, Cout_A1_B22, P_A2_B21, AND_A1_B22, Cout_A1_B21);

    wire AND_A2_B22;
    and and_a2_b22(AND_A2_B22, A[2], B[22]);
    wire P_A2_B22, Cout_A2_B22;
    full_adder add_a2_b22(P_A2_B22, Cout_A2_B22, P_A3_B21, AND_A2_B22, Cout_A2_B21);

    wire AND_A3_B22;
    and and_a3_b22(AND_A3_B22, A[3], B[22]);
    wire P_A3_B22, Cout_A3_B22;
    full_adder add_a3_b22(P_A3_B22, Cout_A3_B22, P_A4_B21, AND_A3_B22, Cout_A3_B21);

    wire AND_A4_B22;
    and and_a4_b22(AND_A4_B22, A[4], B[22]);
    wire P_A4_B22, Cout_A4_B22;
    full_adder add_a4_b22(P_A4_B22, Cout_A4_B22, P_A5_B21, AND_A4_B22, Cout_A4_B21);

    wire AND_A5_B22;
    and and_a5_b22(AND_A5_B22, A[5], B[22]);
    wire P_A5_B22, Cout_A5_B22;
    full_adder add_a5_b22(P_A5_B22, Cout_A5_B22, P_A6_B21, AND_A5_B22, Cout_A5_B21);

    wire AND_A6_B22;
    and and_a6_b22(AND_A6_B22, A[6], B[22]);
    wire P_A6_B22, Cout_A6_B22;
    full_adder add_a6_b22(P_A6_B22, Cout_A6_B22, P_A7_B21, AND_A6_B22, Cout_A6_B21);

    wire AND_A7_B22;
    and and_a7_b22(AND_A7_B22, A[7], B[22]);
    wire P_A7_B22, Cout_A7_B22;
    full_adder add_a7_b22(P_A7_B22, Cout_A7_B22, P_A8_B21, AND_A7_B22, Cout_A7_B21);

    wire AND_A8_B22;
    and and_a8_b22(AND_A8_B22, A[8], B[22]);
    wire P_A8_B22, Cout_A8_B22;
    full_adder add_a8_b22(P_A8_B22, Cout_A8_B22, P_A9_B21, AND_A8_B22, Cout_A8_B21);

    wire AND_A9_B22;
    and and_a9_b22(AND_A9_B22, A[9], B[22]);
    wire P_A9_B22, Cout_A9_B22;
    full_adder add_a9_b22(P_A9_B22, Cout_A9_B22, P_A10_B21, AND_A9_B22, Cout_A9_B21);

    wire AND_A10_B22;
    and and_a10_b22(AND_A10_B22, A[10], B[22]);
    wire P_A10_B22, Cout_A10_B22;
    full_adder add_a10_b22(P_A10_B22, Cout_A10_B22, P_A11_B21, AND_A10_B22, Cout_A10_B21);

    wire AND_A11_B22;
    and and_a11_b22(AND_A11_B22, A[11], B[22]);
    wire P_A11_B22, Cout_A11_B22;
    full_adder add_a11_b22(P_A11_B22, Cout_A11_B22, P_A12_B21, AND_A11_B22, Cout_A11_B21);

    wire AND_A12_B22;
    and and_a12_b22(AND_A12_B22, A[12], B[22]);
    wire P_A12_B22, Cout_A12_B22;
    full_adder add_a12_b22(P_A12_B22, Cout_A12_B22, P_A13_B21, AND_A12_B22, Cout_A12_B21);

    wire AND_A13_B22;
    and and_a13_b22(AND_A13_B22, A[13], B[22]);
    wire P_A13_B22, Cout_A13_B22;
    full_adder add_a13_b22(P_A13_B22, Cout_A13_B22, P_A14_B21, AND_A13_B22, Cout_A13_B21);

    wire AND_A14_B22;
    and and_a14_b22(AND_A14_B22, A[14], B[22]);
    wire P_A14_B22, Cout_A14_B22;
    full_adder add_a14_b22(P_A14_B22, Cout_A14_B22, P_A15_B21, AND_A14_B22, Cout_A14_B21);

    wire AND_A15_B22;
    and and_a15_b22(AND_A15_B22, A[15], B[22]);
    wire P_A15_B22, Cout_A15_B22;
    full_adder add_a15_b22(P_A15_B22, Cout_A15_B22, P_A16_B21, AND_A15_B22, Cout_A15_B21);

    wire AND_A16_B22;
    and and_a16_b22(AND_A16_B22, A[16], B[22]);
    wire P_A16_B22, Cout_A16_B22;
    full_adder add_a16_b22(P_A16_B22, Cout_A16_B22, P_A17_B21, AND_A16_B22, Cout_A16_B21);

    wire AND_A17_B22;
    and and_a17_b22(AND_A17_B22, A[17], B[22]);
    wire P_A17_B22, Cout_A17_B22;
    full_adder add_a17_b22(P_A17_B22, Cout_A17_B22, P_A18_B21, AND_A17_B22, Cout_A17_B21);

    wire AND_A18_B22;
    and and_a18_b22(AND_A18_B22, A[18], B[22]);
    wire P_A18_B22, Cout_A18_B22;
    full_adder add_a18_b22(P_A18_B22, Cout_A18_B22, P_A19_B21, AND_A18_B22, Cout_A18_B21);

    wire AND_A19_B22;
    and and_a19_b22(AND_A19_B22, A[19], B[22]);
    wire P_A19_B22, Cout_A19_B22;
    full_adder add_a19_b22(P_A19_B22, Cout_A19_B22, P_A20_B21, AND_A19_B22, Cout_A19_B21);

    wire AND_A20_B22;
    and and_a20_b22(AND_A20_B22, A[20], B[22]);
    wire P_A20_B22, Cout_A20_B22;
    full_adder add_a20_b22(P_A20_B22, Cout_A20_B22, P_A21_B21, AND_A20_B22, Cout_A20_B21);

    wire AND_A21_B22;
    and and_a21_b22(AND_A21_B22, A[21], B[22]);
    wire P_A21_B22, Cout_A21_B22;
    full_adder add_a21_b22(P_A21_B22, Cout_A21_B22, P_A22_B21, AND_A21_B22, Cout_A21_B21);

    wire AND_A22_B22;
    and and_a22_b22(AND_A22_B22, A[22], B[22]);
    wire P_A22_B22, Cout_A22_B22;
    full_adder add_a22_b22(P_A22_B22, Cout_A22_B22, P_A23_B21, AND_A22_B22, Cout_A22_B21);

    wire AND_A23_B22;
    and and_a23_b22(AND_A23_B22, A[23], B[22]);
    wire P_A23_B22, Cout_A23_B22;
    full_adder add_a23_b22(P_A23_B22, Cout_A23_B22, P_A24_B21, AND_A23_B22, Cout_A23_B21);

    wire AND_A24_B22;
    and and_a24_b22(AND_A24_B22, A[24], B[22]);
    wire P_A24_B22, Cout_A24_B22;
    full_adder add_a24_b22(P_A24_B22, Cout_A24_B22, P_A25_B21, AND_A24_B22, Cout_A24_B21);

    wire AND_A25_B22;
    and and_a25_b22(AND_A25_B22, A[25], B[22]);
    wire P_A25_B22, Cout_A25_B22;
    full_adder add_a25_b22(P_A25_B22, Cout_A25_B22, P_A26_B21, AND_A25_B22, Cout_A25_B21);

    wire AND_A26_B22;
    and and_a26_b22(AND_A26_B22, A[26], B[22]);
    wire P_A26_B22, Cout_A26_B22;
    full_adder add_a26_b22(P_A26_B22, Cout_A26_B22, P_A27_B21, AND_A26_B22, Cout_A26_B21);

    wire AND_A27_B22;
    and and_a27_b22(AND_A27_B22, A[27], B[22]);
    wire P_A27_B22, Cout_A27_B22;
    full_adder add_a27_b22(P_A27_B22, Cout_A27_B22, P_A28_B21, AND_A27_B22, Cout_A27_B21);

    wire AND_A28_B22;
    and and_a28_b22(AND_A28_B22, A[28], B[22]);
    wire P_A28_B22, Cout_A28_B22;
    full_adder add_a28_b22(P_A28_B22, Cout_A28_B22, P_A29_B21, AND_A28_B22, Cout_A28_B21);

    wire AND_A29_B22;
    and and_a29_b22(AND_A29_B22, A[29], B[22]);
    wire P_A29_B22, Cout_A29_B22;
    full_adder add_a29_b22(P_A29_B22, Cout_A29_B22, P_A30_B21, AND_A29_B22, Cout_A29_B21);

    wire AND_A30_B22;
    and and_a30_b22(AND_A30_B22, A[30], B[22]);
    wire P_A30_B22, Cout_A30_B22;
    full_adder add_a30_b22(P_A30_B22, Cout_A30_B22, P_A31_B21, AND_A30_B22, Cout_A30_B21);

    wire AND_A31_B22;
    nand and_a31_b22(AND_A31_B22, A[31], B[22]);
    wire P_A31_B22, Cout_A31_B22;
    half_adder add_a31_b22(P_A31_B22, Cout_A31_B22, AND_A31_B22, Cout_A31_B21);

    wire AND_A0_B23;
    and and_a0_b23(AND_A0_B23, A[0], B[23]);
    wire P_A0_B23, Cout_A0_B23;
    full_adder add_a0_b23(P_A0_B23, Cout_A0_B23, P_A1_B22, AND_A0_B23, Cout_A0_B22);

    wire AND_A1_B23;
    and and_a1_b23(AND_A1_B23, A[1], B[23]);
    wire P_A1_B23, Cout_A1_B23;
    full_adder add_a1_b23(P_A1_B23, Cout_A1_B23, P_A2_B22, AND_A1_B23, Cout_A1_B22);

    wire AND_A2_B23;
    and and_a2_b23(AND_A2_B23, A[2], B[23]);
    wire P_A2_B23, Cout_A2_B23;
    full_adder add_a2_b23(P_A2_B23, Cout_A2_B23, P_A3_B22, AND_A2_B23, Cout_A2_B22);

    wire AND_A3_B23;
    and and_a3_b23(AND_A3_B23, A[3], B[23]);
    wire P_A3_B23, Cout_A3_B23;
    full_adder add_a3_b23(P_A3_B23, Cout_A3_B23, P_A4_B22, AND_A3_B23, Cout_A3_B22);

    wire AND_A4_B23;
    and and_a4_b23(AND_A4_B23, A[4], B[23]);
    wire P_A4_B23, Cout_A4_B23;
    full_adder add_a4_b23(P_A4_B23, Cout_A4_B23, P_A5_B22, AND_A4_B23, Cout_A4_B22);

    wire AND_A5_B23;
    and and_a5_b23(AND_A5_B23, A[5], B[23]);
    wire P_A5_B23, Cout_A5_B23;
    full_adder add_a5_b23(P_A5_B23, Cout_A5_B23, P_A6_B22, AND_A5_B23, Cout_A5_B22);

    wire AND_A6_B23;
    and and_a6_b23(AND_A6_B23, A[6], B[23]);
    wire P_A6_B23, Cout_A6_B23;
    full_adder add_a6_b23(P_A6_B23, Cout_A6_B23, P_A7_B22, AND_A6_B23, Cout_A6_B22);

    wire AND_A7_B23;
    and and_a7_b23(AND_A7_B23, A[7], B[23]);
    wire P_A7_B23, Cout_A7_B23;
    full_adder add_a7_b23(P_A7_B23, Cout_A7_B23, P_A8_B22, AND_A7_B23, Cout_A7_B22);

    wire AND_A8_B23;
    and and_a8_b23(AND_A8_B23, A[8], B[23]);
    wire P_A8_B23, Cout_A8_B23;
    full_adder add_a8_b23(P_A8_B23, Cout_A8_B23, P_A9_B22, AND_A8_B23, Cout_A8_B22);

    wire AND_A9_B23;
    and and_a9_b23(AND_A9_B23, A[9], B[23]);
    wire P_A9_B23, Cout_A9_B23;
    full_adder add_a9_b23(P_A9_B23, Cout_A9_B23, P_A10_B22, AND_A9_B23, Cout_A9_B22);

    wire AND_A10_B23;
    and and_a10_b23(AND_A10_B23, A[10], B[23]);
    wire P_A10_B23, Cout_A10_B23;
    full_adder add_a10_b23(P_A10_B23, Cout_A10_B23, P_A11_B22, AND_A10_B23, Cout_A10_B22);

    wire AND_A11_B23;
    and and_a11_b23(AND_A11_B23, A[11], B[23]);
    wire P_A11_B23, Cout_A11_B23;
    full_adder add_a11_b23(P_A11_B23, Cout_A11_B23, P_A12_B22, AND_A11_B23, Cout_A11_B22);

    wire AND_A12_B23;
    and and_a12_b23(AND_A12_B23, A[12], B[23]);
    wire P_A12_B23, Cout_A12_B23;
    full_adder add_a12_b23(P_A12_B23, Cout_A12_B23, P_A13_B22, AND_A12_B23, Cout_A12_B22);

    wire AND_A13_B23;
    and and_a13_b23(AND_A13_B23, A[13], B[23]);
    wire P_A13_B23, Cout_A13_B23;
    full_adder add_a13_b23(P_A13_B23, Cout_A13_B23, P_A14_B22, AND_A13_B23, Cout_A13_B22);

    wire AND_A14_B23;
    and and_a14_b23(AND_A14_B23, A[14], B[23]);
    wire P_A14_B23, Cout_A14_B23;
    full_adder add_a14_b23(P_A14_B23, Cout_A14_B23, P_A15_B22, AND_A14_B23, Cout_A14_B22);

    wire AND_A15_B23;
    and and_a15_b23(AND_A15_B23, A[15], B[23]);
    wire P_A15_B23, Cout_A15_B23;
    full_adder add_a15_b23(P_A15_B23, Cout_A15_B23, P_A16_B22, AND_A15_B23, Cout_A15_B22);

    wire AND_A16_B23;
    and and_a16_b23(AND_A16_B23, A[16], B[23]);
    wire P_A16_B23, Cout_A16_B23;
    full_adder add_a16_b23(P_A16_B23, Cout_A16_B23, P_A17_B22, AND_A16_B23, Cout_A16_B22);

    wire AND_A17_B23;
    and and_a17_b23(AND_A17_B23, A[17], B[23]);
    wire P_A17_B23, Cout_A17_B23;
    full_adder add_a17_b23(P_A17_B23, Cout_A17_B23, P_A18_B22, AND_A17_B23, Cout_A17_B22);

    wire AND_A18_B23;
    and and_a18_b23(AND_A18_B23, A[18], B[23]);
    wire P_A18_B23, Cout_A18_B23;
    full_adder add_a18_b23(P_A18_B23, Cout_A18_B23, P_A19_B22, AND_A18_B23, Cout_A18_B22);

    wire AND_A19_B23;
    and and_a19_b23(AND_A19_B23, A[19], B[23]);
    wire P_A19_B23, Cout_A19_B23;
    full_adder add_a19_b23(P_A19_B23, Cout_A19_B23, P_A20_B22, AND_A19_B23, Cout_A19_B22);

    wire AND_A20_B23;
    and and_a20_b23(AND_A20_B23, A[20], B[23]);
    wire P_A20_B23, Cout_A20_B23;
    full_adder add_a20_b23(P_A20_B23, Cout_A20_B23, P_A21_B22, AND_A20_B23, Cout_A20_B22);

    wire AND_A21_B23;
    and and_a21_b23(AND_A21_B23, A[21], B[23]);
    wire P_A21_B23, Cout_A21_B23;
    full_adder add_a21_b23(P_A21_B23, Cout_A21_B23, P_A22_B22, AND_A21_B23, Cout_A21_B22);

    wire AND_A22_B23;
    and and_a22_b23(AND_A22_B23, A[22], B[23]);
    wire P_A22_B23, Cout_A22_B23;
    full_adder add_a22_b23(P_A22_B23, Cout_A22_B23, P_A23_B22, AND_A22_B23, Cout_A22_B22);

    wire AND_A23_B23;
    and and_a23_b23(AND_A23_B23, A[23], B[23]);
    wire P_A23_B23, Cout_A23_B23;
    full_adder add_a23_b23(P_A23_B23, Cout_A23_B23, P_A24_B22, AND_A23_B23, Cout_A23_B22);

    wire AND_A24_B23;
    and and_a24_b23(AND_A24_B23, A[24], B[23]);
    wire P_A24_B23, Cout_A24_B23;
    full_adder add_a24_b23(P_A24_B23, Cout_A24_B23, P_A25_B22, AND_A24_B23, Cout_A24_B22);

    wire AND_A25_B23;
    and and_a25_b23(AND_A25_B23, A[25], B[23]);
    wire P_A25_B23, Cout_A25_B23;
    full_adder add_a25_b23(P_A25_B23, Cout_A25_B23, P_A26_B22, AND_A25_B23, Cout_A25_B22);

    wire AND_A26_B23;
    and and_a26_b23(AND_A26_B23, A[26], B[23]);
    wire P_A26_B23, Cout_A26_B23;
    full_adder add_a26_b23(P_A26_B23, Cout_A26_B23, P_A27_B22, AND_A26_B23, Cout_A26_B22);

    wire AND_A27_B23;
    and and_a27_b23(AND_A27_B23, A[27], B[23]);
    wire P_A27_B23, Cout_A27_B23;
    full_adder add_a27_b23(P_A27_B23, Cout_A27_B23, P_A28_B22, AND_A27_B23, Cout_A27_B22);

    wire AND_A28_B23;
    and and_a28_b23(AND_A28_B23, A[28], B[23]);
    wire P_A28_B23, Cout_A28_B23;
    full_adder add_a28_b23(P_A28_B23, Cout_A28_B23, P_A29_B22, AND_A28_B23, Cout_A28_B22);

    wire AND_A29_B23;
    and and_a29_b23(AND_A29_B23, A[29], B[23]);
    wire P_A29_B23, Cout_A29_B23;
    full_adder add_a29_b23(P_A29_B23, Cout_A29_B23, P_A30_B22, AND_A29_B23, Cout_A29_B22);

    wire AND_A30_B23;
    and and_a30_b23(AND_A30_B23, A[30], B[23]);
    wire P_A30_B23, Cout_A30_B23;
    full_adder add_a30_b23(P_A30_B23, Cout_A30_B23, P_A31_B22, AND_A30_B23, Cout_A30_B22);

    wire AND_A31_B23;
    nand and_a31_b23(AND_A31_B23, A[31], B[23]);
    wire P_A31_B23, Cout_A31_B23;
    half_adder add_a31_b23(P_A31_B23, Cout_A31_B23, AND_A31_B23, Cout_A31_B22);

    wire AND_A0_B24;
    and and_a0_b24(AND_A0_B24, A[0], B[24]);
    wire P_A0_B24, Cout_A0_B24;
    full_adder add_a0_b24(P_A0_B24, Cout_A0_B24, P_A1_B23, AND_A0_B24, Cout_A0_B23);

    wire AND_A1_B24;
    and and_a1_b24(AND_A1_B24, A[1], B[24]);
    wire P_A1_B24, Cout_A1_B24;
    full_adder add_a1_b24(P_A1_B24, Cout_A1_B24, P_A2_B23, AND_A1_B24, Cout_A1_B23);

    wire AND_A2_B24;
    and and_a2_b24(AND_A2_B24, A[2], B[24]);
    wire P_A2_B24, Cout_A2_B24;
    full_adder add_a2_b24(P_A2_B24, Cout_A2_B24, P_A3_B23, AND_A2_B24, Cout_A2_B23);

    wire AND_A3_B24;
    and and_a3_b24(AND_A3_B24, A[3], B[24]);
    wire P_A3_B24, Cout_A3_B24;
    full_adder add_a3_b24(P_A3_B24, Cout_A3_B24, P_A4_B23, AND_A3_B24, Cout_A3_B23);

    wire AND_A4_B24;
    and and_a4_b24(AND_A4_B24, A[4], B[24]);
    wire P_A4_B24, Cout_A4_B24;
    full_adder add_a4_b24(P_A4_B24, Cout_A4_B24, P_A5_B23, AND_A4_B24, Cout_A4_B23);

    wire AND_A5_B24;
    and and_a5_b24(AND_A5_B24, A[5], B[24]);
    wire P_A5_B24, Cout_A5_B24;
    full_adder add_a5_b24(P_A5_B24, Cout_A5_B24, P_A6_B23, AND_A5_B24, Cout_A5_B23);

    wire AND_A6_B24;
    and and_a6_b24(AND_A6_B24, A[6], B[24]);
    wire P_A6_B24, Cout_A6_B24;
    full_adder add_a6_b24(P_A6_B24, Cout_A6_B24, P_A7_B23, AND_A6_B24, Cout_A6_B23);

    wire AND_A7_B24;
    and and_a7_b24(AND_A7_B24, A[7], B[24]);
    wire P_A7_B24, Cout_A7_B24;
    full_adder add_a7_b24(P_A7_B24, Cout_A7_B24, P_A8_B23, AND_A7_B24, Cout_A7_B23);

    wire AND_A8_B24;
    and and_a8_b24(AND_A8_B24, A[8], B[24]);
    wire P_A8_B24, Cout_A8_B24;
    full_adder add_a8_b24(P_A8_B24, Cout_A8_B24, P_A9_B23, AND_A8_B24, Cout_A8_B23);

    wire AND_A9_B24;
    and and_a9_b24(AND_A9_B24, A[9], B[24]);
    wire P_A9_B24, Cout_A9_B24;
    full_adder add_a9_b24(P_A9_B24, Cout_A9_B24, P_A10_B23, AND_A9_B24, Cout_A9_B23);

    wire AND_A10_B24;
    and and_a10_b24(AND_A10_B24, A[10], B[24]);
    wire P_A10_B24, Cout_A10_B24;
    full_adder add_a10_b24(P_A10_B24, Cout_A10_B24, P_A11_B23, AND_A10_B24, Cout_A10_B23);

    wire AND_A11_B24;
    and and_a11_b24(AND_A11_B24, A[11], B[24]);
    wire P_A11_B24, Cout_A11_B24;
    full_adder add_a11_b24(P_A11_B24, Cout_A11_B24, P_A12_B23, AND_A11_B24, Cout_A11_B23);

    wire AND_A12_B24;
    and and_a12_b24(AND_A12_B24, A[12], B[24]);
    wire P_A12_B24, Cout_A12_B24;
    full_adder add_a12_b24(P_A12_B24, Cout_A12_B24, P_A13_B23, AND_A12_B24, Cout_A12_B23);

    wire AND_A13_B24;
    and and_a13_b24(AND_A13_B24, A[13], B[24]);
    wire P_A13_B24, Cout_A13_B24;
    full_adder add_a13_b24(P_A13_B24, Cout_A13_B24, P_A14_B23, AND_A13_B24, Cout_A13_B23);

    wire AND_A14_B24;
    and and_a14_b24(AND_A14_B24, A[14], B[24]);
    wire P_A14_B24, Cout_A14_B24;
    full_adder add_a14_b24(P_A14_B24, Cout_A14_B24, P_A15_B23, AND_A14_B24, Cout_A14_B23);

    wire AND_A15_B24;
    and and_a15_b24(AND_A15_B24, A[15], B[24]);
    wire P_A15_B24, Cout_A15_B24;
    full_adder add_a15_b24(P_A15_B24, Cout_A15_B24, P_A16_B23, AND_A15_B24, Cout_A15_B23);

    wire AND_A16_B24;
    and and_a16_b24(AND_A16_B24, A[16], B[24]);
    wire P_A16_B24, Cout_A16_B24;
    full_adder add_a16_b24(P_A16_B24, Cout_A16_B24, P_A17_B23, AND_A16_B24, Cout_A16_B23);

    wire AND_A17_B24;
    and and_a17_b24(AND_A17_B24, A[17], B[24]);
    wire P_A17_B24, Cout_A17_B24;
    full_adder add_a17_b24(P_A17_B24, Cout_A17_B24, P_A18_B23, AND_A17_B24, Cout_A17_B23);

    wire AND_A18_B24;
    and and_a18_b24(AND_A18_B24, A[18], B[24]);
    wire P_A18_B24, Cout_A18_B24;
    full_adder add_a18_b24(P_A18_B24, Cout_A18_B24, P_A19_B23, AND_A18_B24, Cout_A18_B23);

    wire AND_A19_B24;
    and and_a19_b24(AND_A19_B24, A[19], B[24]);
    wire P_A19_B24, Cout_A19_B24;
    full_adder add_a19_b24(P_A19_B24, Cout_A19_B24, P_A20_B23, AND_A19_B24, Cout_A19_B23);

    wire AND_A20_B24;
    and and_a20_b24(AND_A20_B24, A[20], B[24]);
    wire P_A20_B24, Cout_A20_B24;
    full_adder add_a20_b24(P_A20_B24, Cout_A20_B24, P_A21_B23, AND_A20_B24, Cout_A20_B23);

    wire AND_A21_B24;
    and and_a21_b24(AND_A21_B24, A[21], B[24]);
    wire P_A21_B24, Cout_A21_B24;
    full_adder add_a21_b24(P_A21_B24, Cout_A21_B24, P_A22_B23, AND_A21_B24, Cout_A21_B23);

    wire AND_A22_B24;
    and and_a22_b24(AND_A22_B24, A[22], B[24]);
    wire P_A22_B24, Cout_A22_B24;
    full_adder add_a22_b24(P_A22_B24, Cout_A22_B24, P_A23_B23, AND_A22_B24, Cout_A22_B23);

    wire AND_A23_B24;
    and and_a23_b24(AND_A23_B24, A[23], B[24]);
    wire P_A23_B24, Cout_A23_B24;
    full_adder add_a23_b24(P_A23_B24, Cout_A23_B24, P_A24_B23, AND_A23_B24, Cout_A23_B23);

    wire AND_A24_B24;
    and and_a24_b24(AND_A24_B24, A[24], B[24]);
    wire P_A24_B24, Cout_A24_B24;
    full_adder add_a24_b24(P_A24_B24, Cout_A24_B24, P_A25_B23, AND_A24_B24, Cout_A24_B23);

    wire AND_A25_B24;
    and and_a25_b24(AND_A25_B24, A[25], B[24]);
    wire P_A25_B24, Cout_A25_B24;
    full_adder add_a25_b24(P_A25_B24, Cout_A25_B24, P_A26_B23, AND_A25_B24, Cout_A25_B23);

    wire AND_A26_B24;
    and and_a26_b24(AND_A26_B24, A[26], B[24]);
    wire P_A26_B24, Cout_A26_B24;
    full_adder add_a26_b24(P_A26_B24, Cout_A26_B24, P_A27_B23, AND_A26_B24, Cout_A26_B23);

    wire AND_A27_B24;
    and and_a27_b24(AND_A27_B24, A[27], B[24]);
    wire P_A27_B24, Cout_A27_B24;
    full_adder add_a27_b24(P_A27_B24, Cout_A27_B24, P_A28_B23, AND_A27_B24, Cout_A27_B23);

    wire AND_A28_B24;
    and and_a28_b24(AND_A28_B24, A[28], B[24]);
    wire P_A28_B24, Cout_A28_B24;
    full_adder add_a28_b24(P_A28_B24, Cout_A28_B24, P_A29_B23, AND_A28_B24, Cout_A28_B23);

    wire AND_A29_B24;
    and and_a29_b24(AND_A29_B24, A[29], B[24]);
    wire P_A29_B24, Cout_A29_B24;
    full_adder add_a29_b24(P_A29_B24, Cout_A29_B24, P_A30_B23, AND_A29_B24, Cout_A29_B23);

    wire AND_A30_B24;
    and and_a30_b24(AND_A30_B24, A[30], B[24]);
    wire P_A30_B24, Cout_A30_B24;
    full_adder add_a30_b24(P_A30_B24, Cout_A30_B24, P_A31_B23, AND_A30_B24, Cout_A30_B23);

    wire AND_A31_B24;
    nand and_a31_b24(AND_A31_B24, A[31], B[24]);
    wire P_A31_B24, Cout_A31_B24;
    half_adder add_a31_b24(P_A31_B24, Cout_A31_B24, AND_A31_B24, Cout_A31_B23);

    wire AND_A0_B25;
    and and_a0_b25(AND_A0_B25, A[0], B[25]);
    wire P_A0_B25, Cout_A0_B25;
    full_adder add_a0_b25(P_A0_B25, Cout_A0_B25, P_A1_B24, AND_A0_B25, Cout_A0_B24);

    wire AND_A1_B25;
    and and_a1_b25(AND_A1_B25, A[1], B[25]);
    wire P_A1_B25, Cout_A1_B25;
    full_adder add_a1_b25(P_A1_B25, Cout_A1_B25, P_A2_B24, AND_A1_B25, Cout_A1_B24);

    wire AND_A2_B25;
    and and_a2_b25(AND_A2_B25, A[2], B[25]);
    wire P_A2_B25, Cout_A2_B25;
    full_adder add_a2_b25(P_A2_B25, Cout_A2_B25, P_A3_B24, AND_A2_B25, Cout_A2_B24);

    wire AND_A3_B25;
    and and_a3_b25(AND_A3_B25, A[3], B[25]);
    wire P_A3_B25, Cout_A3_B25;
    full_adder add_a3_b25(P_A3_B25, Cout_A3_B25, P_A4_B24, AND_A3_B25, Cout_A3_B24);

    wire AND_A4_B25;
    and and_a4_b25(AND_A4_B25, A[4], B[25]);
    wire P_A4_B25, Cout_A4_B25;
    full_adder add_a4_b25(P_A4_B25, Cout_A4_B25, P_A5_B24, AND_A4_B25, Cout_A4_B24);

    wire AND_A5_B25;
    and and_a5_b25(AND_A5_B25, A[5], B[25]);
    wire P_A5_B25, Cout_A5_B25;
    full_adder add_a5_b25(P_A5_B25, Cout_A5_B25, P_A6_B24, AND_A5_B25, Cout_A5_B24);

    wire AND_A6_B25;
    and and_a6_b25(AND_A6_B25, A[6], B[25]);
    wire P_A6_B25, Cout_A6_B25;
    full_adder add_a6_b25(P_A6_B25, Cout_A6_B25, P_A7_B24, AND_A6_B25, Cout_A6_B24);

    wire AND_A7_B25;
    and and_a7_b25(AND_A7_B25, A[7], B[25]);
    wire P_A7_B25, Cout_A7_B25;
    full_adder add_a7_b25(P_A7_B25, Cout_A7_B25, P_A8_B24, AND_A7_B25, Cout_A7_B24);

    wire AND_A8_B25;
    and and_a8_b25(AND_A8_B25, A[8], B[25]);
    wire P_A8_B25, Cout_A8_B25;
    full_adder add_a8_b25(P_A8_B25, Cout_A8_B25, P_A9_B24, AND_A8_B25, Cout_A8_B24);

    wire AND_A9_B25;
    and and_a9_b25(AND_A9_B25, A[9], B[25]);
    wire P_A9_B25, Cout_A9_B25;
    full_adder add_a9_b25(P_A9_B25, Cout_A9_B25, P_A10_B24, AND_A9_B25, Cout_A9_B24);

    wire AND_A10_B25;
    and and_a10_b25(AND_A10_B25, A[10], B[25]);
    wire P_A10_B25, Cout_A10_B25;
    full_adder add_a10_b25(P_A10_B25, Cout_A10_B25, P_A11_B24, AND_A10_B25, Cout_A10_B24);

    wire AND_A11_B25;
    and and_a11_b25(AND_A11_B25, A[11], B[25]);
    wire P_A11_B25, Cout_A11_B25;
    full_adder add_a11_b25(P_A11_B25, Cout_A11_B25, P_A12_B24, AND_A11_B25, Cout_A11_B24);

    wire AND_A12_B25;
    and and_a12_b25(AND_A12_B25, A[12], B[25]);
    wire P_A12_B25, Cout_A12_B25;
    full_adder add_a12_b25(P_A12_B25, Cout_A12_B25, P_A13_B24, AND_A12_B25, Cout_A12_B24);

    wire AND_A13_B25;
    and and_a13_b25(AND_A13_B25, A[13], B[25]);
    wire P_A13_B25, Cout_A13_B25;
    full_adder add_a13_b25(P_A13_B25, Cout_A13_B25, P_A14_B24, AND_A13_B25, Cout_A13_B24);

    wire AND_A14_B25;
    and and_a14_b25(AND_A14_B25, A[14], B[25]);
    wire P_A14_B25, Cout_A14_B25;
    full_adder add_a14_b25(P_A14_B25, Cout_A14_B25, P_A15_B24, AND_A14_B25, Cout_A14_B24);

    wire AND_A15_B25;
    and and_a15_b25(AND_A15_B25, A[15], B[25]);
    wire P_A15_B25, Cout_A15_B25;
    full_adder add_a15_b25(P_A15_B25, Cout_A15_B25, P_A16_B24, AND_A15_B25, Cout_A15_B24);

    wire AND_A16_B25;
    and and_a16_b25(AND_A16_B25, A[16], B[25]);
    wire P_A16_B25, Cout_A16_B25;
    full_adder add_a16_b25(P_A16_B25, Cout_A16_B25, P_A17_B24, AND_A16_B25, Cout_A16_B24);

    wire AND_A17_B25;
    and and_a17_b25(AND_A17_B25, A[17], B[25]);
    wire P_A17_B25, Cout_A17_B25;
    full_adder add_a17_b25(P_A17_B25, Cout_A17_B25, P_A18_B24, AND_A17_B25, Cout_A17_B24);

    wire AND_A18_B25;
    and and_a18_b25(AND_A18_B25, A[18], B[25]);
    wire P_A18_B25, Cout_A18_B25;
    full_adder add_a18_b25(P_A18_B25, Cout_A18_B25, P_A19_B24, AND_A18_B25, Cout_A18_B24);

    wire AND_A19_B25;
    and and_a19_b25(AND_A19_B25, A[19], B[25]);
    wire P_A19_B25, Cout_A19_B25;
    full_adder add_a19_b25(P_A19_B25, Cout_A19_B25, P_A20_B24, AND_A19_B25, Cout_A19_B24);

    wire AND_A20_B25;
    and and_a20_b25(AND_A20_B25, A[20], B[25]);
    wire P_A20_B25, Cout_A20_B25;
    full_adder add_a20_b25(P_A20_B25, Cout_A20_B25, P_A21_B24, AND_A20_B25, Cout_A20_B24);

    wire AND_A21_B25;
    and and_a21_b25(AND_A21_B25, A[21], B[25]);
    wire P_A21_B25, Cout_A21_B25;
    full_adder add_a21_b25(P_A21_B25, Cout_A21_B25, P_A22_B24, AND_A21_B25, Cout_A21_B24);

    wire AND_A22_B25;
    and and_a22_b25(AND_A22_B25, A[22], B[25]);
    wire P_A22_B25, Cout_A22_B25;
    full_adder add_a22_b25(P_A22_B25, Cout_A22_B25, P_A23_B24, AND_A22_B25, Cout_A22_B24);

    wire AND_A23_B25;
    and and_a23_b25(AND_A23_B25, A[23], B[25]);
    wire P_A23_B25, Cout_A23_B25;
    full_adder add_a23_b25(P_A23_B25, Cout_A23_B25, P_A24_B24, AND_A23_B25, Cout_A23_B24);

    wire AND_A24_B25;
    and and_a24_b25(AND_A24_B25, A[24], B[25]);
    wire P_A24_B25, Cout_A24_B25;
    full_adder add_a24_b25(P_A24_B25, Cout_A24_B25, P_A25_B24, AND_A24_B25, Cout_A24_B24);

    wire AND_A25_B25;
    and and_a25_b25(AND_A25_B25, A[25], B[25]);
    wire P_A25_B25, Cout_A25_B25;
    full_adder add_a25_b25(P_A25_B25, Cout_A25_B25, P_A26_B24, AND_A25_B25, Cout_A25_B24);

    wire AND_A26_B25;
    and and_a26_b25(AND_A26_B25, A[26], B[25]);
    wire P_A26_B25, Cout_A26_B25;
    full_adder add_a26_b25(P_A26_B25, Cout_A26_B25, P_A27_B24, AND_A26_B25, Cout_A26_B24);

    wire AND_A27_B25;
    and and_a27_b25(AND_A27_B25, A[27], B[25]);
    wire P_A27_B25, Cout_A27_B25;
    full_adder add_a27_b25(P_A27_B25, Cout_A27_B25, P_A28_B24, AND_A27_B25, Cout_A27_B24);

    wire AND_A28_B25;
    and and_a28_b25(AND_A28_B25, A[28], B[25]);
    wire P_A28_B25, Cout_A28_B25;
    full_adder add_a28_b25(P_A28_B25, Cout_A28_B25, P_A29_B24, AND_A28_B25, Cout_A28_B24);

    wire AND_A29_B25;
    and and_a29_b25(AND_A29_B25, A[29], B[25]);
    wire P_A29_B25, Cout_A29_B25;
    full_adder add_a29_b25(P_A29_B25, Cout_A29_B25, P_A30_B24, AND_A29_B25, Cout_A29_B24);

    wire AND_A30_B25;
    and and_a30_b25(AND_A30_B25, A[30], B[25]);
    wire P_A30_B25, Cout_A30_B25;
    full_adder add_a30_b25(P_A30_B25, Cout_A30_B25, P_A31_B24, AND_A30_B25, Cout_A30_B24);

    wire AND_A31_B25;
    nand and_a31_b25(AND_A31_B25, A[31], B[25]);
    wire P_A31_B25, Cout_A31_B25;
    half_adder add_a31_b25(P_A31_B25, Cout_A31_B25, AND_A31_B25, Cout_A31_B24);

    wire AND_A0_B26;
    and and_a0_b26(AND_A0_B26, A[0], B[26]);
    wire P_A0_B26, Cout_A0_B26;
    full_adder add_a0_b26(P_A0_B26, Cout_A0_B26, P_A1_B25, AND_A0_B26, Cout_A0_B25);

    wire AND_A1_B26;
    and and_a1_b26(AND_A1_B26, A[1], B[26]);
    wire P_A1_B26, Cout_A1_B26;
    full_adder add_a1_b26(P_A1_B26, Cout_A1_B26, P_A2_B25, AND_A1_B26, Cout_A1_B25);

    wire AND_A2_B26;
    and and_a2_b26(AND_A2_B26, A[2], B[26]);
    wire P_A2_B26, Cout_A2_B26;
    full_adder add_a2_b26(P_A2_B26, Cout_A2_B26, P_A3_B25, AND_A2_B26, Cout_A2_B25);

    wire AND_A3_B26;
    and and_a3_b26(AND_A3_B26, A[3], B[26]);
    wire P_A3_B26, Cout_A3_B26;
    full_adder add_a3_b26(P_A3_B26, Cout_A3_B26, P_A4_B25, AND_A3_B26, Cout_A3_B25);

    wire AND_A4_B26;
    and and_a4_b26(AND_A4_B26, A[4], B[26]);
    wire P_A4_B26, Cout_A4_B26;
    full_adder add_a4_b26(P_A4_B26, Cout_A4_B26, P_A5_B25, AND_A4_B26, Cout_A4_B25);

    wire AND_A5_B26;
    and and_a5_b26(AND_A5_B26, A[5], B[26]);
    wire P_A5_B26, Cout_A5_B26;
    full_adder add_a5_b26(P_A5_B26, Cout_A5_B26, P_A6_B25, AND_A5_B26, Cout_A5_B25);

    wire AND_A6_B26;
    and and_a6_b26(AND_A6_B26, A[6], B[26]);
    wire P_A6_B26, Cout_A6_B26;
    full_adder add_a6_b26(P_A6_B26, Cout_A6_B26, P_A7_B25, AND_A6_B26, Cout_A6_B25);

    wire AND_A7_B26;
    and and_a7_b26(AND_A7_B26, A[7], B[26]);
    wire P_A7_B26, Cout_A7_B26;
    full_adder add_a7_b26(P_A7_B26, Cout_A7_B26, P_A8_B25, AND_A7_B26, Cout_A7_B25);

    wire AND_A8_B26;
    and and_a8_b26(AND_A8_B26, A[8], B[26]);
    wire P_A8_B26, Cout_A8_B26;
    full_adder add_a8_b26(P_A8_B26, Cout_A8_B26, P_A9_B25, AND_A8_B26, Cout_A8_B25);

    wire AND_A9_B26;
    and and_a9_b26(AND_A9_B26, A[9], B[26]);
    wire P_A9_B26, Cout_A9_B26;
    full_adder add_a9_b26(P_A9_B26, Cout_A9_B26, P_A10_B25, AND_A9_B26, Cout_A9_B25);

    wire AND_A10_B26;
    and and_a10_b26(AND_A10_B26, A[10], B[26]);
    wire P_A10_B26, Cout_A10_B26;
    full_adder add_a10_b26(P_A10_B26, Cout_A10_B26, P_A11_B25, AND_A10_B26, Cout_A10_B25);

    wire AND_A11_B26;
    and and_a11_b26(AND_A11_B26, A[11], B[26]);
    wire P_A11_B26, Cout_A11_B26;
    full_adder add_a11_b26(P_A11_B26, Cout_A11_B26, P_A12_B25, AND_A11_B26, Cout_A11_B25);

    wire AND_A12_B26;
    and and_a12_b26(AND_A12_B26, A[12], B[26]);
    wire P_A12_B26, Cout_A12_B26;
    full_adder add_a12_b26(P_A12_B26, Cout_A12_B26, P_A13_B25, AND_A12_B26, Cout_A12_B25);

    wire AND_A13_B26;
    and and_a13_b26(AND_A13_B26, A[13], B[26]);
    wire P_A13_B26, Cout_A13_B26;
    full_adder add_a13_b26(P_A13_B26, Cout_A13_B26, P_A14_B25, AND_A13_B26, Cout_A13_B25);

    wire AND_A14_B26;
    and and_a14_b26(AND_A14_B26, A[14], B[26]);
    wire P_A14_B26, Cout_A14_B26;
    full_adder add_a14_b26(P_A14_B26, Cout_A14_B26, P_A15_B25, AND_A14_B26, Cout_A14_B25);

    wire AND_A15_B26;
    and and_a15_b26(AND_A15_B26, A[15], B[26]);
    wire P_A15_B26, Cout_A15_B26;
    full_adder add_a15_b26(P_A15_B26, Cout_A15_B26, P_A16_B25, AND_A15_B26, Cout_A15_B25);

    wire AND_A16_B26;
    and and_a16_b26(AND_A16_B26, A[16], B[26]);
    wire P_A16_B26, Cout_A16_B26;
    full_adder add_a16_b26(P_A16_B26, Cout_A16_B26, P_A17_B25, AND_A16_B26, Cout_A16_B25);

    wire AND_A17_B26;
    and and_a17_b26(AND_A17_B26, A[17], B[26]);
    wire P_A17_B26, Cout_A17_B26;
    full_adder add_a17_b26(P_A17_B26, Cout_A17_B26, P_A18_B25, AND_A17_B26, Cout_A17_B25);

    wire AND_A18_B26;
    and and_a18_b26(AND_A18_B26, A[18], B[26]);
    wire P_A18_B26, Cout_A18_B26;
    full_adder add_a18_b26(P_A18_B26, Cout_A18_B26, P_A19_B25, AND_A18_B26, Cout_A18_B25);

    wire AND_A19_B26;
    and and_a19_b26(AND_A19_B26, A[19], B[26]);
    wire P_A19_B26, Cout_A19_B26;
    full_adder add_a19_b26(P_A19_B26, Cout_A19_B26, P_A20_B25, AND_A19_B26, Cout_A19_B25);

    wire AND_A20_B26;
    and and_a20_b26(AND_A20_B26, A[20], B[26]);
    wire P_A20_B26, Cout_A20_B26;
    full_adder add_a20_b26(P_A20_B26, Cout_A20_B26, P_A21_B25, AND_A20_B26, Cout_A20_B25);

    wire AND_A21_B26;
    and and_a21_b26(AND_A21_B26, A[21], B[26]);
    wire P_A21_B26, Cout_A21_B26;
    full_adder add_a21_b26(P_A21_B26, Cout_A21_B26, P_A22_B25, AND_A21_B26, Cout_A21_B25);

    wire AND_A22_B26;
    and and_a22_b26(AND_A22_B26, A[22], B[26]);
    wire P_A22_B26, Cout_A22_B26;
    full_adder add_a22_b26(P_A22_B26, Cout_A22_B26, P_A23_B25, AND_A22_B26, Cout_A22_B25);

    wire AND_A23_B26;
    and and_a23_b26(AND_A23_B26, A[23], B[26]);
    wire P_A23_B26, Cout_A23_B26;
    full_adder add_a23_b26(P_A23_B26, Cout_A23_B26, P_A24_B25, AND_A23_B26, Cout_A23_B25);

    wire AND_A24_B26;
    and and_a24_b26(AND_A24_B26, A[24], B[26]);
    wire P_A24_B26, Cout_A24_B26;
    full_adder add_a24_b26(P_A24_B26, Cout_A24_B26, P_A25_B25, AND_A24_B26, Cout_A24_B25);

    wire AND_A25_B26;
    and and_a25_b26(AND_A25_B26, A[25], B[26]);
    wire P_A25_B26, Cout_A25_B26;
    full_adder add_a25_b26(P_A25_B26, Cout_A25_B26, P_A26_B25, AND_A25_B26, Cout_A25_B25);

    wire AND_A26_B26;
    and and_a26_b26(AND_A26_B26, A[26], B[26]);
    wire P_A26_B26, Cout_A26_B26;
    full_adder add_a26_b26(P_A26_B26, Cout_A26_B26, P_A27_B25, AND_A26_B26, Cout_A26_B25);

    wire AND_A27_B26;
    and and_a27_b26(AND_A27_B26, A[27], B[26]);
    wire P_A27_B26, Cout_A27_B26;
    full_adder add_a27_b26(P_A27_B26, Cout_A27_B26, P_A28_B25, AND_A27_B26, Cout_A27_B25);

    wire AND_A28_B26;
    and and_a28_b26(AND_A28_B26, A[28], B[26]);
    wire P_A28_B26, Cout_A28_B26;
    full_adder add_a28_b26(P_A28_B26, Cout_A28_B26, P_A29_B25, AND_A28_B26, Cout_A28_B25);

    wire AND_A29_B26;
    and and_a29_b26(AND_A29_B26, A[29], B[26]);
    wire P_A29_B26, Cout_A29_B26;
    full_adder add_a29_b26(P_A29_B26, Cout_A29_B26, P_A30_B25, AND_A29_B26, Cout_A29_B25);

    wire AND_A30_B26;
    and and_a30_b26(AND_A30_B26, A[30], B[26]);
    wire P_A30_B26, Cout_A30_B26;
    full_adder add_a30_b26(P_A30_B26, Cout_A30_B26, P_A31_B25, AND_A30_B26, Cout_A30_B25);

    wire AND_A31_B26;
    nand and_a31_b26(AND_A31_B26, A[31], B[26]);
    wire P_A31_B26, Cout_A31_B26;
    half_adder add_a31_b26(P_A31_B26, Cout_A31_B26, AND_A31_B26, Cout_A31_B25);

    wire AND_A0_B27;
    and and_a0_b27(AND_A0_B27, A[0], B[27]);
    wire P_A0_B27, Cout_A0_B27;
    full_adder add_a0_b27(P_A0_B27, Cout_A0_B27, P_A1_B26, AND_A0_B27, Cout_A0_B26);

    wire AND_A1_B27;
    and and_a1_b27(AND_A1_B27, A[1], B[27]);
    wire P_A1_B27, Cout_A1_B27;
    full_adder add_a1_b27(P_A1_B27, Cout_A1_B27, P_A2_B26, AND_A1_B27, Cout_A1_B26);

    wire AND_A2_B27;
    and and_a2_b27(AND_A2_B27, A[2], B[27]);
    wire P_A2_B27, Cout_A2_B27;
    full_adder add_a2_b27(P_A2_B27, Cout_A2_B27, P_A3_B26, AND_A2_B27, Cout_A2_B26);

    wire AND_A3_B27;
    and and_a3_b27(AND_A3_B27, A[3], B[27]);
    wire P_A3_B27, Cout_A3_B27;
    full_adder add_a3_b27(P_A3_B27, Cout_A3_B27, P_A4_B26, AND_A3_B27, Cout_A3_B26);

    wire AND_A4_B27;
    and and_a4_b27(AND_A4_B27, A[4], B[27]);
    wire P_A4_B27, Cout_A4_B27;
    full_adder add_a4_b27(P_A4_B27, Cout_A4_B27, P_A5_B26, AND_A4_B27, Cout_A4_B26);

    wire AND_A5_B27;
    and and_a5_b27(AND_A5_B27, A[5], B[27]);
    wire P_A5_B27, Cout_A5_B27;
    full_adder add_a5_b27(P_A5_B27, Cout_A5_B27, P_A6_B26, AND_A5_B27, Cout_A5_B26);

    wire AND_A6_B27;
    and and_a6_b27(AND_A6_B27, A[6], B[27]);
    wire P_A6_B27, Cout_A6_B27;
    full_adder add_a6_b27(P_A6_B27, Cout_A6_B27, P_A7_B26, AND_A6_B27, Cout_A6_B26);

    wire AND_A7_B27;
    and and_a7_b27(AND_A7_B27, A[7], B[27]);
    wire P_A7_B27, Cout_A7_B27;
    full_adder add_a7_b27(P_A7_B27, Cout_A7_B27, P_A8_B26, AND_A7_B27, Cout_A7_B26);

    wire AND_A8_B27;
    and and_a8_b27(AND_A8_B27, A[8], B[27]);
    wire P_A8_B27, Cout_A8_B27;
    full_adder add_a8_b27(P_A8_B27, Cout_A8_B27, P_A9_B26, AND_A8_B27, Cout_A8_B26);

    wire AND_A9_B27;
    and and_a9_b27(AND_A9_B27, A[9], B[27]);
    wire P_A9_B27, Cout_A9_B27;
    full_adder add_a9_b27(P_A9_B27, Cout_A9_B27, P_A10_B26, AND_A9_B27, Cout_A9_B26);

    wire AND_A10_B27;
    and and_a10_b27(AND_A10_B27, A[10], B[27]);
    wire P_A10_B27, Cout_A10_B27;
    full_adder add_a10_b27(P_A10_B27, Cout_A10_B27, P_A11_B26, AND_A10_B27, Cout_A10_B26);

    wire AND_A11_B27;
    and and_a11_b27(AND_A11_B27, A[11], B[27]);
    wire P_A11_B27, Cout_A11_B27;
    full_adder add_a11_b27(P_A11_B27, Cout_A11_B27, P_A12_B26, AND_A11_B27, Cout_A11_B26);

    wire AND_A12_B27;
    and and_a12_b27(AND_A12_B27, A[12], B[27]);
    wire P_A12_B27, Cout_A12_B27;
    full_adder add_a12_b27(P_A12_B27, Cout_A12_B27, P_A13_B26, AND_A12_B27, Cout_A12_B26);

    wire AND_A13_B27;
    and and_a13_b27(AND_A13_B27, A[13], B[27]);
    wire P_A13_B27, Cout_A13_B27;
    full_adder add_a13_b27(P_A13_B27, Cout_A13_B27, P_A14_B26, AND_A13_B27, Cout_A13_B26);

    wire AND_A14_B27;
    and and_a14_b27(AND_A14_B27, A[14], B[27]);
    wire P_A14_B27, Cout_A14_B27;
    full_adder add_a14_b27(P_A14_B27, Cout_A14_B27, P_A15_B26, AND_A14_B27, Cout_A14_B26);

    wire AND_A15_B27;
    and and_a15_b27(AND_A15_B27, A[15], B[27]);
    wire P_A15_B27, Cout_A15_B27;
    full_adder add_a15_b27(P_A15_B27, Cout_A15_B27, P_A16_B26, AND_A15_B27, Cout_A15_B26);

    wire AND_A16_B27;
    and and_a16_b27(AND_A16_B27, A[16], B[27]);
    wire P_A16_B27, Cout_A16_B27;
    full_adder add_a16_b27(P_A16_B27, Cout_A16_B27, P_A17_B26, AND_A16_B27, Cout_A16_B26);

    wire AND_A17_B27;
    and and_a17_b27(AND_A17_B27, A[17], B[27]);
    wire P_A17_B27, Cout_A17_B27;
    full_adder add_a17_b27(P_A17_B27, Cout_A17_B27, P_A18_B26, AND_A17_B27, Cout_A17_B26);

    wire AND_A18_B27;
    and and_a18_b27(AND_A18_B27, A[18], B[27]);
    wire P_A18_B27, Cout_A18_B27;
    full_adder add_a18_b27(P_A18_B27, Cout_A18_B27, P_A19_B26, AND_A18_B27, Cout_A18_B26);

    wire AND_A19_B27;
    and and_a19_b27(AND_A19_B27, A[19], B[27]);
    wire P_A19_B27, Cout_A19_B27;
    full_adder add_a19_b27(P_A19_B27, Cout_A19_B27, P_A20_B26, AND_A19_B27, Cout_A19_B26);

    wire AND_A20_B27;
    and and_a20_b27(AND_A20_B27, A[20], B[27]);
    wire P_A20_B27, Cout_A20_B27;
    full_adder add_a20_b27(P_A20_B27, Cout_A20_B27, P_A21_B26, AND_A20_B27, Cout_A20_B26);

    wire AND_A21_B27;
    and and_a21_b27(AND_A21_B27, A[21], B[27]);
    wire P_A21_B27, Cout_A21_B27;
    full_adder add_a21_b27(P_A21_B27, Cout_A21_B27, P_A22_B26, AND_A21_B27, Cout_A21_B26);

    wire AND_A22_B27;
    and and_a22_b27(AND_A22_B27, A[22], B[27]);
    wire P_A22_B27, Cout_A22_B27;
    full_adder add_a22_b27(P_A22_B27, Cout_A22_B27, P_A23_B26, AND_A22_B27, Cout_A22_B26);

    wire AND_A23_B27;
    and and_a23_b27(AND_A23_B27, A[23], B[27]);
    wire P_A23_B27, Cout_A23_B27;
    full_adder add_a23_b27(P_A23_B27, Cout_A23_B27, P_A24_B26, AND_A23_B27, Cout_A23_B26);

    wire AND_A24_B27;
    and and_a24_b27(AND_A24_B27, A[24], B[27]);
    wire P_A24_B27, Cout_A24_B27;
    full_adder add_a24_b27(P_A24_B27, Cout_A24_B27, P_A25_B26, AND_A24_B27, Cout_A24_B26);

    wire AND_A25_B27;
    and and_a25_b27(AND_A25_B27, A[25], B[27]);
    wire P_A25_B27, Cout_A25_B27;
    full_adder add_a25_b27(P_A25_B27, Cout_A25_B27, P_A26_B26, AND_A25_B27, Cout_A25_B26);

    wire AND_A26_B27;
    and and_a26_b27(AND_A26_B27, A[26], B[27]);
    wire P_A26_B27, Cout_A26_B27;
    full_adder add_a26_b27(P_A26_B27, Cout_A26_B27, P_A27_B26, AND_A26_B27, Cout_A26_B26);

    wire AND_A27_B27;
    and and_a27_b27(AND_A27_B27, A[27], B[27]);
    wire P_A27_B27, Cout_A27_B27;
    full_adder add_a27_b27(P_A27_B27, Cout_A27_B27, P_A28_B26, AND_A27_B27, Cout_A27_B26);

    wire AND_A28_B27;
    and and_a28_b27(AND_A28_B27, A[28], B[27]);
    wire P_A28_B27, Cout_A28_B27;
    full_adder add_a28_b27(P_A28_B27, Cout_A28_B27, P_A29_B26, AND_A28_B27, Cout_A28_B26);

    wire AND_A29_B27;
    and and_a29_b27(AND_A29_B27, A[29], B[27]);
    wire P_A29_B27, Cout_A29_B27;
    full_adder add_a29_b27(P_A29_B27, Cout_A29_B27, P_A30_B26, AND_A29_B27, Cout_A29_B26);

    wire AND_A30_B27;
    and and_a30_b27(AND_A30_B27, A[30], B[27]);
    wire P_A30_B27, Cout_A30_B27;
    full_adder add_a30_b27(P_A30_B27, Cout_A30_B27, P_A31_B26, AND_A30_B27, Cout_A30_B26);

    wire AND_A31_B27;
    nand and_a31_b27(AND_A31_B27, A[31], B[27]);
    wire P_A31_B27, Cout_A31_B27;
    half_adder add_a31_b27(P_A31_B27, Cout_A31_B27, AND_A31_B27, Cout_A31_B26);

    wire AND_A0_B28;
    and and_a0_b28(AND_A0_B28, A[0], B[28]);
    wire P_A0_B28, Cout_A0_B28;
    full_adder add_a0_b28(P_A0_B28, Cout_A0_B28, P_A1_B27, AND_A0_B28, Cout_A0_B27);

    wire AND_A1_B28;
    and and_a1_b28(AND_A1_B28, A[1], B[28]);
    wire P_A1_B28, Cout_A1_B28;
    full_adder add_a1_b28(P_A1_B28, Cout_A1_B28, P_A2_B27, AND_A1_B28, Cout_A1_B27);

    wire AND_A2_B28;
    and and_a2_b28(AND_A2_B28, A[2], B[28]);
    wire P_A2_B28, Cout_A2_B28;
    full_adder add_a2_b28(P_A2_B28, Cout_A2_B28, P_A3_B27, AND_A2_B28, Cout_A2_B27);

    wire AND_A3_B28;
    and and_a3_b28(AND_A3_B28, A[3], B[28]);
    wire P_A3_B28, Cout_A3_B28;
    full_adder add_a3_b28(P_A3_B28, Cout_A3_B28, P_A4_B27, AND_A3_B28, Cout_A3_B27);

    wire AND_A4_B28;
    and and_a4_b28(AND_A4_B28, A[4], B[28]);
    wire P_A4_B28, Cout_A4_B28;
    full_adder add_a4_b28(P_A4_B28, Cout_A4_B28, P_A5_B27, AND_A4_B28, Cout_A4_B27);

    wire AND_A5_B28;
    and and_a5_b28(AND_A5_B28, A[5], B[28]);
    wire P_A5_B28, Cout_A5_B28;
    full_adder add_a5_b28(P_A5_B28, Cout_A5_B28, P_A6_B27, AND_A5_B28, Cout_A5_B27);

    wire AND_A6_B28;
    and and_a6_b28(AND_A6_B28, A[6], B[28]);
    wire P_A6_B28, Cout_A6_B28;
    full_adder add_a6_b28(P_A6_B28, Cout_A6_B28, P_A7_B27, AND_A6_B28, Cout_A6_B27);

    wire AND_A7_B28;
    and and_a7_b28(AND_A7_B28, A[7], B[28]);
    wire P_A7_B28, Cout_A7_B28;
    full_adder add_a7_b28(P_A7_B28, Cout_A7_B28, P_A8_B27, AND_A7_B28, Cout_A7_B27);

    wire AND_A8_B28;
    and and_a8_b28(AND_A8_B28, A[8], B[28]);
    wire P_A8_B28, Cout_A8_B28;
    full_adder add_a8_b28(P_A8_B28, Cout_A8_B28, P_A9_B27, AND_A8_B28, Cout_A8_B27);

    wire AND_A9_B28;
    and and_a9_b28(AND_A9_B28, A[9], B[28]);
    wire P_A9_B28, Cout_A9_B28;
    full_adder add_a9_b28(P_A9_B28, Cout_A9_B28, P_A10_B27, AND_A9_B28, Cout_A9_B27);

    wire AND_A10_B28;
    and and_a10_b28(AND_A10_B28, A[10], B[28]);
    wire P_A10_B28, Cout_A10_B28;
    full_adder add_a10_b28(P_A10_B28, Cout_A10_B28, P_A11_B27, AND_A10_B28, Cout_A10_B27);

    wire AND_A11_B28;
    and and_a11_b28(AND_A11_B28, A[11], B[28]);
    wire P_A11_B28, Cout_A11_B28;
    full_adder add_a11_b28(P_A11_B28, Cout_A11_B28, P_A12_B27, AND_A11_B28, Cout_A11_B27);

    wire AND_A12_B28;
    and and_a12_b28(AND_A12_B28, A[12], B[28]);
    wire P_A12_B28, Cout_A12_B28;
    full_adder add_a12_b28(P_A12_B28, Cout_A12_B28, P_A13_B27, AND_A12_B28, Cout_A12_B27);

    wire AND_A13_B28;
    and and_a13_b28(AND_A13_B28, A[13], B[28]);
    wire P_A13_B28, Cout_A13_B28;
    full_adder add_a13_b28(P_A13_B28, Cout_A13_B28, P_A14_B27, AND_A13_B28, Cout_A13_B27);

    wire AND_A14_B28;
    and and_a14_b28(AND_A14_B28, A[14], B[28]);
    wire P_A14_B28, Cout_A14_B28;
    full_adder add_a14_b28(P_A14_B28, Cout_A14_B28, P_A15_B27, AND_A14_B28, Cout_A14_B27);

    wire AND_A15_B28;
    and and_a15_b28(AND_A15_B28, A[15], B[28]);
    wire P_A15_B28, Cout_A15_B28;
    full_adder add_a15_b28(P_A15_B28, Cout_A15_B28, P_A16_B27, AND_A15_B28, Cout_A15_B27);

    wire AND_A16_B28;
    and and_a16_b28(AND_A16_B28, A[16], B[28]);
    wire P_A16_B28, Cout_A16_B28;
    full_adder add_a16_b28(P_A16_B28, Cout_A16_B28, P_A17_B27, AND_A16_B28, Cout_A16_B27);

    wire AND_A17_B28;
    and and_a17_b28(AND_A17_B28, A[17], B[28]);
    wire P_A17_B28, Cout_A17_B28;
    full_adder add_a17_b28(P_A17_B28, Cout_A17_B28, P_A18_B27, AND_A17_B28, Cout_A17_B27);

    wire AND_A18_B28;
    and and_a18_b28(AND_A18_B28, A[18], B[28]);
    wire P_A18_B28, Cout_A18_B28;
    full_adder add_a18_b28(P_A18_B28, Cout_A18_B28, P_A19_B27, AND_A18_B28, Cout_A18_B27);

    wire AND_A19_B28;
    and and_a19_b28(AND_A19_B28, A[19], B[28]);
    wire P_A19_B28, Cout_A19_B28;
    full_adder add_a19_b28(P_A19_B28, Cout_A19_B28, P_A20_B27, AND_A19_B28, Cout_A19_B27);

    wire AND_A20_B28;
    and and_a20_b28(AND_A20_B28, A[20], B[28]);
    wire P_A20_B28, Cout_A20_B28;
    full_adder add_a20_b28(P_A20_B28, Cout_A20_B28, P_A21_B27, AND_A20_B28, Cout_A20_B27);

    wire AND_A21_B28;
    and and_a21_b28(AND_A21_B28, A[21], B[28]);
    wire P_A21_B28, Cout_A21_B28;
    full_adder add_a21_b28(P_A21_B28, Cout_A21_B28, P_A22_B27, AND_A21_B28, Cout_A21_B27);

    wire AND_A22_B28;
    and and_a22_b28(AND_A22_B28, A[22], B[28]);
    wire P_A22_B28, Cout_A22_B28;
    full_adder add_a22_b28(P_A22_B28, Cout_A22_B28, P_A23_B27, AND_A22_B28, Cout_A22_B27);

    wire AND_A23_B28;
    and and_a23_b28(AND_A23_B28, A[23], B[28]);
    wire P_A23_B28, Cout_A23_B28;
    full_adder add_a23_b28(P_A23_B28, Cout_A23_B28, P_A24_B27, AND_A23_B28, Cout_A23_B27);

    wire AND_A24_B28;
    and and_a24_b28(AND_A24_B28, A[24], B[28]);
    wire P_A24_B28, Cout_A24_B28;
    full_adder add_a24_b28(P_A24_B28, Cout_A24_B28, P_A25_B27, AND_A24_B28, Cout_A24_B27);

    wire AND_A25_B28;
    and and_a25_b28(AND_A25_B28, A[25], B[28]);
    wire P_A25_B28, Cout_A25_B28;
    full_adder add_a25_b28(P_A25_B28, Cout_A25_B28, P_A26_B27, AND_A25_B28, Cout_A25_B27);

    wire AND_A26_B28;
    and and_a26_b28(AND_A26_B28, A[26], B[28]);
    wire P_A26_B28, Cout_A26_B28;
    full_adder add_a26_b28(P_A26_B28, Cout_A26_B28, P_A27_B27, AND_A26_B28, Cout_A26_B27);

    wire AND_A27_B28;
    and and_a27_b28(AND_A27_B28, A[27], B[28]);
    wire P_A27_B28, Cout_A27_B28;
    full_adder add_a27_b28(P_A27_B28, Cout_A27_B28, P_A28_B27, AND_A27_B28, Cout_A27_B27);

    wire AND_A28_B28;
    and and_a28_b28(AND_A28_B28, A[28], B[28]);
    wire P_A28_B28, Cout_A28_B28;
    full_adder add_a28_b28(P_A28_B28, Cout_A28_B28, P_A29_B27, AND_A28_B28, Cout_A28_B27);

    wire AND_A29_B28;
    and and_a29_b28(AND_A29_B28, A[29], B[28]);
    wire P_A29_B28, Cout_A29_B28;
    full_adder add_a29_b28(P_A29_B28, Cout_A29_B28, P_A30_B27, AND_A29_B28, Cout_A29_B27);

    wire AND_A30_B28;
    and and_a30_b28(AND_A30_B28, A[30], B[28]);
    wire P_A30_B28, Cout_A30_B28;
    full_adder add_a30_b28(P_A30_B28, Cout_A30_B28, P_A31_B27, AND_A30_B28, Cout_A30_B27);

    wire AND_A31_B28;
    nand and_a31_b28(AND_A31_B28, A[31], B[28]);
    wire P_A31_B28, Cout_A31_B28;
    half_adder add_a31_b28(P_A31_B28, Cout_A31_B28, AND_A31_B28, Cout_A31_B27);

    wire AND_A0_B29;
    and and_a0_b29(AND_A0_B29, A[0], B[29]);
    wire P_A0_B29, Cout_A0_B29;
    full_adder add_a0_b29(P_A0_B29, Cout_A0_B29, P_A1_B28, AND_A0_B29, Cout_A0_B28);

    wire AND_A1_B29;
    and and_a1_b29(AND_A1_B29, A[1], B[29]);
    wire P_A1_B29, Cout_A1_B29;
    full_adder add_a1_b29(P_A1_B29, Cout_A1_B29, P_A2_B28, AND_A1_B29, Cout_A1_B28);

    wire AND_A2_B29;
    and and_a2_b29(AND_A2_B29, A[2], B[29]);
    wire P_A2_B29, Cout_A2_B29;
    full_adder add_a2_b29(P_A2_B29, Cout_A2_B29, P_A3_B28, AND_A2_B29, Cout_A2_B28);

    wire AND_A3_B29;
    and and_a3_b29(AND_A3_B29, A[3], B[29]);
    wire P_A3_B29, Cout_A3_B29;
    full_adder add_a3_b29(P_A3_B29, Cout_A3_B29, P_A4_B28, AND_A3_B29, Cout_A3_B28);

    wire AND_A4_B29;
    and and_a4_b29(AND_A4_B29, A[4], B[29]);
    wire P_A4_B29, Cout_A4_B29;
    full_adder add_a4_b29(P_A4_B29, Cout_A4_B29, P_A5_B28, AND_A4_B29, Cout_A4_B28);

    wire AND_A5_B29;
    and and_a5_b29(AND_A5_B29, A[5], B[29]);
    wire P_A5_B29, Cout_A5_B29;
    full_adder add_a5_b29(P_A5_B29, Cout_A5_B29, P_A6_B28, AND_A5_B29, Cout_A5_B28);

    wire AND_A6_B29;
    and and_a6_b29(AND_A6_B29, A[6], B[29]);
    wire P_A6_B29, Cout_A6_B29;
    full_adder add_a6_b29(P_A6_B29, Cout_A6_B29, P_A7_B28, AND_A6_B29, Cout_A6_B28);

    wire AND_A7_B29;
    and and_a7_b29(AND_A7_B29, A[7], B[29]);
    wire P_A7_B29, Cout_A7_B29;
    full_adder add_a7_b29(P_A7_B29, Cout_A7_B29, P_A8_B28, AND_A7_B29, Cout_A7_B28);

    wire AND_A8_B29;
    and and_a8_b29(AND_A8_B29, A[8], B[29]);
    wire P_A8_B29, Cout_A8_B29;
    full_adder add_a8_b29(P_A8_B29, Cout_A8_B29, P_A9_B28, AND_A8_B29, Cout_A8_B28);

    wire AND_A9_B29;
    and and_a9_b29(AND_A9_B29, A[9], B[29]);
    wire P_A9_B29, Cout_A9_B29;
    full_adder add_a9_b29(P_A9_B29, Cout_A9_B29, P_A10_B28, AND_A9_B29, Cout_A9_B28);

    wire AND_A10_B29;
    and and_a10_b29(AND_A10_B29, A[10], B[29]);
    wire P_A10_B29, Cout_A10_B29;
    full_adder add_a10_b29(P_A10_B29, Cout_A10_B29, P_A11_B28, AND_A10_B29, Cout_A10_B28);

    wire AND_A11_B29;
    and and_a11_b29(AND_A11_B29, A[11], B[29]);
    wire P_A11_B29, Cout_A11_B29;
    full_adder add_a11_b29(P_A11_B29, Cout_A11_B29, P_A12_B28, AND_A11_B29, Cout_A11_B28);

    wire AND_A12_B29;
    and and_a12_b29(AND_A12_B29, A[12], B[29]);
    wire P_A12_B29, Cout_A12_B29;
    full_adder add_a12_b29(P_A12_B29, Cout_A12_B29, P_A13_B28, AND_A12_B29, Cout_A12_B28);

    wire AND_A13_B29;
    and and_a13_b29(AND_A13_B29, A[13], B[29]);
    wire P_A13_B29, Cout_A13_B29;
    full_adder add_a13_b29(P_A13_B29, Cout_A13_B29, P_A14_B28, AND_A13_B29, Cout_A13_B28);

    wire AND_A14_B29;
    and and_a14_b29(AND_A14_B29, A[14], B[29]);
    wire P_A14_B29, Cout_A14_B29;
    full_adder add_a14_b29(P_A14_B29, Cout_A14_B29, P_A15_B28, AND_A14_B29, Cout_A14_B28);

    wire AND_A15_B29;
    and and_a15_b29(AND_A15_B29, A[15], B[29]);
    wire P_A15_B29, Cout_A15_B29;
    full_adder add_a15_b29(P_A15_B29, Cout_A15_B29, P_A16_B28, AND_A15_B29, Cout_A15_B28);

    wire AND_A16_B29;
    and and_a16_b29(AND_A16_B29, A[16], B[29]);
    wire P_A16_B29, Cout_A16_B29;
    full_adder add_a16_b29(P_A16_B29, Cout_A16_B29, P_A17_B28, AND_A16_B29, Cout_A16_B28);

    wire AND_A17_B29;
    and and_a17_b29(AND_A17_B29, A[17], B[29]);
    wire P_A17_B29, Cout_A17_B29;
    full_adder add_a17_b29(P_A17_B29, Cout_A17_B29, P_A18_B28, AND_A17_B29, Cout_A17_B28);

    wire AND_A18_B29;
    and and_a18_b29(AND_A18_B29, A[18], B[29]);
    wire P_A18_B29, Cout_A18_B29;
    full_adder add_a18_b29(P_A18_B29, Cout_A18_B29, P_A19_B28, AND_A18_B29, Cout_A18_B28);

    wire AND_A19_B29;
    and and_a19_b29(AND_A19_B29, A[19], B[29]);
    wire P_A19_B29, Cout_A19_B29;
    full_adder add_a19_b29(P_A19_B29, Cout_A19_B29, P_A20_B28, AND_A19_B29, Cout_A19_B28);

    wire AND_A20_B29;
    and and_a20_b29(AND_A20_B29, A[20], B[29]);
    wire P_A20_B29, Cout_A20_B29;
    full_adder add_a20_b29(P_A20_B29, Cout_A20_B29, P_A21_B28, AND_A20_B29, Cout_A20_B28);

    wire AND_A21_B29;
    and and_a21_b29(AND_A21_B29, A[21], B[29]);
    wire P_A21_B29, Cout_A21_B29;
    full_adder add_a21_b29(P_A21_B29, Cout_A21_B29, P_A22_B28, AND_A21_B29, Cout_A21_B28);

    wire AND_A22_B29;
    and and_a22_b29(AND_A22_B29, A[22], B[29]);
    wire P_A22_B29, Cout_A22_B29;
    full_adder add_a22_b29(P_A22_B29, Cout_A22_B29, P_A23_B28, AND_A22_B29, Cout_A22_B28);

    wire AND_A23_B29;
    and and_a23_b29(AND_A23_B29, A[23], B[29]);
    wire P_A23_B29, Cout_A23_B29;
    full_adder add_a23_b29(P_A23_B29, Cout_A23_B29, P_A24_B28, AND_A23_B29, Cout_A23_B28);

    wire AND_A24_B29;
    and and_a24_b29(AND_A24_B29, A[24], B[29]);
    wire P_A24_B29, Cout_A24_B29;
    full_adder add_a24_b29(P_A24_B29, Cout_A24_B29, P_A25_B28, AND_A24_B29, Cout_A24_B28);

    wire AND_A25_B29;
    and and_a25_b29(AND_A25_B29, A[25], B[29]);
    wire P_A25_B29, Cout_A25_B29;
    full_adder add_a25_b29(P_A25_B29, Cout_A25_B29, P_A26_B28, AND_A25_B29, Cout_A25_B28);

    wire AND_A26_B29;
    and and_a26_b29(AND_A26_B29, A[26], B[29]);
    wire P_A26_B29, Cout_A26_B29;
    full_adder add_a26_b29(P_A26_B29, Cout_A26_B29, P_A27_B28, AND_A26_B29, Cout_A26_B28);

    wire AND_A27_B29;
    and and_a27_b29(AND_A27_B29, A[27], B[29]);
    wire P_A27_B29, Cout_A27_B29;
    full_adder add_a27_b29(P_A27_B29, Cout_A27_B29, P_A28_B28, AND_A27_B29, Cout_A27_B28);

    wire AND_A28_B29;
    and and_a28_b29(AND_A28_B29, A[28], B[29]);
    wire P_A28_B29, Cout_A28_B29;
    full_adder add_a28_b29(P_A28_B29, Cout_A28_B29, P_A29_B28, AND_A28_B29, Cout_A28_B28);

    wire AND_A29_B29;
    and and_a29_b29(AND_A29_B29, A[29], B[29]);
    wire P_A29_B29, Cout_A29_B29;
    full_adder add_a29_b29(P_A29_B29, Cout_A29_B29, P_A30_B28, AND_A29_B29, Cout_A29_B28);

    wire AND_A30_B29;
    and and_a30_b29(AND_A30_B29, A[30], B[29]);
    wire P_A30_B29, Cout_A30_B29;
    full_adder add_a30_b29(P_A30_B29, Cout_A30_B29, P_A31_B28, AND_A30_B29, Cout_A30_B28);

    wire AND_A31_B29;
    nand and_a31_b29(AND_A31_B29, A[31], B[29]);
    wire P_A31_B29, Cout_A31_B29;
    half_adder add_a31_b29(P_A31_B29, Cout_A31_B29, AND_A31_B29, Cout_A31_B28);

    wire AND_A0_B30;
    and and_a0_b30(AND_A0_B30, A[0], B[30]);
    wire P_A0_B30, Cout_A0_B30;
    full_adder add_a0_b30(P_A0_B30, Cout_A0_B30, P_A1_B29, AND_A0_B30, Cout_A0_B29);

    wire AND_A1_B30;
    and and_a1_b30(AND_A1_B30, A[1], B[30]);
    wire P_A1_B30, Cout_A1_B30;
    full_adder add_a1_b30(P_A1_B30, Cout_A1_B30, P_A2_B29, AND_A1_B30, Cout_A1_B29);

    wire AND_A2_B30;
    and and_a2_b30(AND_A2_B30, A[2], B[30]);
    wire P_A2_B30, Cout_A2_B30;
    full_adder add_a2_b30(P_A2_B30, Cout_A2_B30, P_A3_B29, AND_A2_B30, Cout_A2_B29);

    wire AND_A3_B30;
    and and_a3_b30(AND_A3_B30, A[3], B[30]);
    wire P_A3_B30, Cout_A3_B30;
    full_adder add_a3_b30(P_A3_B30, Cout_A3_B30, P_A4_B29, AND_A3_B30, Cout_A3_B29);

    wire AND_A4_B30;
    and and_a4_b30(AND_A4_B30, A[4], B[30]);
    wire P_A4_B30, Cout_A4_B30;
    full_adder add_a4_b30(P_A4_B30, Cout_A4_B30, P_A5_B29, AND_A4_B30, Cout_A4_B29);

    wire AND_A5_B30;
    and and_a5_b30(AND_A5_B30, A[5], B[30]);
    wire P_A5_B30, Cout_A5_B30;
    full_adder add_a5_b30(P_A5_B30, Cout_A5_B30, P_A6_B29, AND_A5_B30, Cout_A5_B29);

    wire AND_A6_B30;
    and and_a6_b30(AND_A6_B30, A[6], B[30]);
    wire P_A6_B30, Cout_A6_B30;
    full_adder add_a6_b30(P_A6_B30, Cout_A6_B30, P_A7_B29, AND_A6_B30, Cout_A6_B29);

    wire AND_A7_B30;
    and and_a7_b30(AND_A7_B30, A[7], B[30]);
    wire P_A7_B30, Cout_A7_B30;
    full_adder add_a7_b30(P_A7_B30, Cout_A7_B30, P_A8_B29, AND_A7_B30, Cout_A7_B29);

    wire AND_A8_B30;
    and and_a8_b30(AND_A8_B30, A[8], B[30]);
    wire P_A8_B30, Cout_A8_B30;
    full_adder add_a8_b30(P_A8_B30, Cout_A8_B30, P_A9_B29, AND_A8_B30, Cout_A8_B29);

    wire AND_A9_B30;
    and and_a9_b30(AND_A9_B30, A[9], B[30]);
    wire P_A9_B30, Cout_A9_B30;
    full_adder add_a9_b30(P_A9_B30, Cout_A9_B30, P_A10_B29, AND_A9_B30, Cout_A9_B29);

    wire AND_A10_B30;
    and and_a10_b30(AND_A10_B30, A[10], B[30]);
    wire P_A10_B30, Cout_A10_B30;
    full_adder add_a10_b30(P_A10_B30, Cout_A10_B30, P_A11_B29, AND_A10_B30, Cout_A10_B29);

    wire AND_A11_B30;
    and and_a11_b30(AND_A11_B30, A[11], B[30]);
    wire P_A11_B30, Cout_A11_B30;
    full_adder add_a11_b30(P_A11_B30, Cout_A11_B30, P_A12_B29, AND_A11_B30, Cout_A11_B29);

    wire AND_A12_B30;
    and and_a12_b30(AND_A12_B30, A[12], B[30]);
    wire P_A12_B30, Cout_A12_B30;
    full_adder add_a12_b30(P_A12_B30, Cout_A12_B30, P_A13_B29, AND_A12_B30, Cout_A12_B29);

    wire AND_A13_B30;
    and and_a13_b30(AND_A13_B30, A[13], B[30]);
    wire P_A13_B30, Cout_A13_B30;
    full_adder add_a13_b30(P_A13_B30, Cout_A13_B30, P_A14_B29, AND_A13_B30, Cout_A13_B29);

    wire AND_A14_B30;
    and and_a14_b30(AND_A14_B30, A[14], B[30]);
    wire P_A14_B30, Cout_A14_B30;
    full_adder add_a14_b30(P_A14_B30, Cout_A14_B30, P_A15_B29, AND_A14_B30, Cout_A14_B29);

    wire AND_A15_B30;
    and and_a15_b30(AND_A15_B30, A[15], B[30]);
    wire P_A15_B30, Cout_A15_B30;
    full_adder add_a15_b30(P_A15_B30, Cout_A15_B30, P_A16_B29, AND_A15_B30, Cout_A15_B29);

    wire AND_A16_B30;
    and and_a16_b30(AND_A16_B30, A[16], B[30]);
    wire P_A16_B30, Cout_A16_B30;
    full_adder add_a16_b30(P_A16_B30, Cout_A16_B30, P_A17_B29, AND_A16_B30, Cout_A16_B29);

    wire AND_A17_B30;
    and and_a17_b30(AND_A17_B30, A[17], B[30]);
    wire P_A17_B30, Cout_A17_B30;
    full_adder add_a17_b30(P_A17_B30, Cout_A17_B30, P_A18_B29, AND_A17_B30, Cout_A17_B29);

    wire AND_A18_B30;
    and and_a18_b30(AND_A18_B30, A[18], B[30]);
    wire P_A18_B30, Cout_A18_B30;
    full_adder add_a18_b30(P_A18_B30, Cout_A18_B30, P_A19_B29, AND_A18_B30, Cout_A18_B29);

    wire AND_A19_B30;
    and and_a19_b30(AND_A19_B30, A[19], B[30]);
    wire P_A19_B30, Cout_A19_B30;
    full_adder add_a19_b30(P_A19_B30, Cout_A19_B30, P_A20_B29, AND_A19_B30, Cout_A19_B29);

    wire AND_A20_B30;
    and and_a20_b30(AND_A20_B30, A[20], B[30]);
    wire P_A20_B30, Cout_A20_B30;
    full_adder add_a20_b30(P_A20_B30, Cout_A20_B30, P_A21_B29, AND_A20_B30, Cout_A20_B29);

    wire AND_A21_B30;
    and and_a21_b30(AND_A21_B30, A[21], B[30]);
    wire P_A21_B30, Cout_A21_B30;
    full_adder add_a21_b30(P_A21_B30, Cout_A21_B30, P_A22_B29, AND_A21_B30, Cout_A21_B29);

    wire AND_A22_B30;
    and and_a22_b30(AND_A22_B30, A[22], B[30]);
    wire P_A22_B30, Cout_A22_B30;
    full_adder add_a22_b30(P_A22_B30, Cout_A22_B30, P_A23_B29, AND_A22_B30, Cout_A22_B29);

    wire AND_A23_B30;
    and and_a23_b30(AND_A23_B30, A[23], B[30]);
    wire P_A23_B30, Cout_A23_B30;
    full_adder add_a23_b30(P_A23_B30, Cout_A23_B30, P_A24_B29, AND_A23_B30, Cout_A23_B29);

    wire AND_A24_B30;
    and and_a24_b30(AND_A24_B30, A[24], B[30]);
    wire P_A24_B30, Cout_A24_B30;
    full_adder add_a24_b30(P_A24_B30, Cout_A24_B30, P_A25_B29, AND_A24_B30, Cout_A24_B29);

    wire AND_A25_B30;
    and and_a25_b30(AND_A25_B30, A[25], B[30]);
    wire P_A25_B30, Cout_A25_B30;
    full_adder add_a25_b30(P_A25_B30, Cout_A25_B30, P_A26_B29, AND_A25_B30, Cout_A25_B29);

    wire AND_A26_B30;
    and and_a26_b30(AND_A26_B30, A[26], B[30]);
    wire P_A26_B30, Cout_A26_B30;
    full_adder add_a26_b30(P_A26_B30, Cout_A26_B30, P_A27_B29, AND_A26_B30, Cout_A26_B29);

    wire AND_A27_B30;
    and and_a27_b30(AND_A27_B30, A[27], B[30]);
    wire P_A27_B30, Cout_A27_B30;
    full_adder add_a27_b30(P_A27_B30, Cout_A27_B30, P_A28_B29, AND_A27_B30, Cout_A27_B29);

    wire AND_A28_B30;
    and and_a28_b30(AND_A28_B30, A[28], B[30]);
    wire P_A28_B30, Cout_A28_B30;
    full_adder add_a28_b30(P_A28_B30, Cout_A28_B30, P_A29_B29, AND_A28_B30, Cout_A28_B29);

    wire AND_A29_B30;
    and and_a29_b30(AND_A29_B30, A[29], B[30]);
    wire P_A29_B30, Cout_A29_B30;
    full_adder add_a29_b30(P_A29_B30, Cout_A29_B30, P_A30_B29, AND_A29_B30, Cout_A29_B29);

    wire AND_A30_B30;
    and and_a30_b30(AND_A30_B30, A[30], B[30]);
    wire P_A30_B30, Cout_A30_B30;
    full_adder add_a30_b30(P_A30_B30, Cout_A30_B30, P_A31_B29, AND_A30_B30, Cout_A30_B29);

    wire AND_A31_B30;
    nand and_a31_b30(AND_A31_B30, A[31], B[30]);
    wire P_A31_B30, Cout_A31_B30;
    half_adder add_a31_b30(P_A31_B30, Cout_A31_B30, AND_A31_B30, Cout_A31_B29);

    wire AND_A0_B31;
    nand and_a0_b31(AND_A0_B31, A[0], B[31]);
    wire P_A0_B31, Cout_A0_B31;
    full_adder add_a0_b31(P_A0_B31, Cout_A0_B31, P_A1_B30, AND_A0_B31, Cout_A0_B30);

    wire AND_A1_B31;
    nand and_a1_b31(AND_A1_B31, A[1], B[31]);
    wire P_A1_B31, Cout_A1_B31;
    full_adder add_a1_b31(P_A1_B31, Cout_A1_B31, P_A2_B30, AND_A1_B31, Cout_A1_B30);

    wire AND_A2_B31;
    nand and_a2_b31(AND_A2_B31, A[2], B[31]);
    wire P_A2_B31, Cout_A2_B31;
    full_adder add_a2_b31(P_A2_B31, Cout_A2_B31, P_A3_B30, AND_A2_B31, Cout_A2_B30);

    wire AND_A3_B31;
    nand and_a3_b31(AND_A3_B31, A[3], B[31]);
    wire P_A3_B31, Cout_A3_B31;
    full_adder add_a3_b31(P_A3_B31, Cout_A3_B31, P_A4_B30, AND_A3_B31, Cout_A3_B30);

    wire AND_A4_B31;
    nand and_a4_b31(AND_A4_B31, A[4], B[31]);
    wire P_A4_B31, Cout_A4_B31;
    full_adder add_a4_b31(P_A4_B31, Cout_A4_B31, P_A5_B30, AND_A4_B31, Cout_A4_B30);

    wire AND_A5_B31;
    nand and_a5_b31(AND_A5_B31, A[5], B[31]);
    wire P_A5_B31, Cout_A5_B31;
    full_adder add_a5_b31(P_A5_B31, Cout_A5_B31, P_A6_B30, AND_A5_B31, Cout_A5_B30);

    wire AND_A6_B31;
    nand and_a6_b31(AND_A6_B31, A[6], B[31]);
    wire P_A6_B31, Cout_A6_B31;
    full_adder add_a6_b31(P_A6_B31, Cout_A6_B31, P_A7_B30, AND_A6_B31, Cout_A6_B30);

    wire AND_A7_B31;
    nand and_a7_b31(AND_A7_B31, A[7], B[31]);
    wire P_A7_B31, Cout_A7_B31;
    full_adder add_a7_b31(P_A7_B31, Cout_A7_B31, P_A8_B30, AND_A7_B31, Cout_A7_B30);

    wire AND_A8_B31;
    nand and_a8_b31(AND_A8_B31, A[8], B[31]);
    wire P_A8_B31, Cout_A8_B31;
    full_adder add_a8_b31(P_A8_B31, Cout_A8_B31, P_A9_B30, AND_A8_B31, Cout_A8_B30);

    wire AND_A9_B31;
    nand and_a9_b31(AND_A9_B31, A[9], B[31]);
    wire P_A9_B31, Cout_A9_B31;
    full_adder add_a9_b31(P_A9_B31, Cout_A9_B31, P_A10_B30, AND_A9_B31, Cout_A9_B30);

    wire AND_A10_B31;
    nand and_a10_b31(AND_A10_B31, A[10], B[31]);
    wire P_A10_B31, Cout_A10_B31;
    full_adder add_a10_b31(P_A10_B31, Cout_A10_B31, P_A11_B30, AND_A10_B31, Cout_A10_B30);

    wire AND_A11_B31;
    nand and_a11_b31(AND_A11_B31, A[11], B[31]);
    wire P_A11_B31, Cout_A11_B31;
    full_adder add_a11_b31(P_A11_B31, Cout_A11_B31, P_A12_B30, AND_A11_B31, Cout_A11_B30);

    wire AND_A12_B31;
    nand and_a12_b31(AND_A12_B31, A[12], B[31]);
    wire P_A12_B31, Cout_A12_B31;
    full_adder add_a12_b31(P_A12_B31, Cout_A12_B31, P_A13_B30, AND_A12_B31, Cout_A12_B30);

    wire AND_A13_B31;
    nand and_a13_b31(AND_A13_B31, A[13], B[31]);
    wire P_A13_B31, Cout_A13_B31;
    full_adder add_a13_b31(P_A13_B31, Cout_A13_B31, P_A14_B30, AND_A13_B31, Cout_A13_B30);

    wire AND_A14_B31;
    nand and_a14_b31(AND_A14_B31, A[14], B[31]);
    wire P_A14_B31, Cout_A14_B31;
    full_adder add_a14_b31(P_A14_B31, Cout_A14_B31, P_A15_B30, AND_A14_B31, Cout_A14_B30);

    wire AND_A15_B31;
    nand and_a15_b31(AND_A15_B31, A[15], B[31]);
    wire P_A15_B31, Cout_A15_B31;
    full_adder add_a15_b31(P_A15_B31, Cout_A15_B31, P_A16_B30, AND_A15_B31, Cout_A15_B30);

    wire AND_A16_B31;
    nand and_a16_b31(AND_A16_B31, A[16], B[31]);
    wire P_A16_B31, Cout_A16_B31;
    full_adder add_a16_b31(P_A16_B31, Cout_A16_B31, P_A17_B30, AND_A16_B31, Cout_A16_B30);

    wire AND_A17_B31;
    nand and_a17_b31(AND_A17_B31, A[17], B[31]);
    wire P_A17_B31, Cout_A17_B31;
    full_adder add_a17_b31(P_A17_B31, Cout_A17_B31, P_A18_B30, AND_A17_B31, Cout_A17_B30);

    wire AND_A18_B31;
    nand and_a18_b31(AND_A18_B31, A[18], B[31]);
    wire P_A18_B31, Cout_A18_B31;
    full_adder add_a18_b31(P_A18_B31, Cout_A18_B31, P_A19_B30, AND_A18_B31, Cout_A18_B30);

    wire AND_A19_B31;
    nand and_a19_b31(AND_A19_B31, A[19], B[31]);
    wire P_A19_B31, Cout_A19_B31;
    full_adder add_a19_b31(P_A19_B31, Cout_A19_B31, P_A20_B30, AND_A19_B31, Cout_A19_B30);

    wire AND_A20_B31;
    nand and_a20_b31(AND_A20_B31, A[20], B[31]);
    wire P_A20_B31, Cout_A20_B31;
    full_adder add_a20_b31(P_A20_B31, Cout_A20_B31, P_A21_B30, AND_A20_B31, Cout_A20_B30);

    wire AND_A21_B31;
    nand and_a21_b31(AND_A21_B31, A[21], B[31]);
    wire P_A21_B31, Cout_A21_B31;
    full_adder add_a21_b31(P_A21_B31, Cout_A21_B31, P_A22_B30, AND_A21_B31, Cout_A21_B30);

    wire AND_A22_B31;
    nand and_a22_b31(AND_A22_B31, A[22], B[31]);
    wire P_A22_B31, Cout_A22_B31;
    full_adder add_a22_b31(P_A22_B31, Cout_A22_B31, P_A23_B30, AND_A22_B31, Cout_A22_B30);

    wire AND_A23_B31;
    nand and_a23_b31(AND_A23_B31, A[23], B[31]);
    wire P_A23_B31, Cout_A23_B31;
    full_adder add_a23_b31(P_A23_B31, Cout_A23_B31, P_A24_B30, AND_A23_B31, Cout_A23_B30);

    wire AND_A24_B31;
    nand and_a24_b31(AND_A24_B31, A[24], B[31]);
    wire P_A24_B31, Cout_A24_B31;
    full_adder add_a24_b31(P_A24_B31, Cout_A24_B31, P_A25_B30, AND_A24_B31, Cout_A24_B30);

    wire AND_A25_B31;
    nand and_a25_b31(AND_A25_B31, A[25], B[31]);
    wire P_A25_B31, Cout_A25_B31;
    full_adder add_a25_b31(P_A25_B31, Cout_A25_B31, P_A26_B30, AND_A25_B31, Cout_A25_B30);

    wire AND_A26_B31;
    nand and_a26_b31(AND_A26_B31, A[26], B[31]);
    wire P_A26_B31, Cout_A26_B31;
    full_adder add_a26_b31(P_A26_B31, Cout_A26_B31, P_A27_B30, AND_A26_B31, Cout_A26_B30);

    wire AND_A27_B31;
    nand and_a27_b31(AND_A27_B31, A[27], B[31]);
    wire P_A27_B31, Cout_A27_B31;
    full_adder add_a27_b31(P_A27_B31, Cout_A27_B31, P_A28_B30, AND_A27_B31, Cout_A27_B30);

    wire AND_A28_B31;
    nand and_a28_b31(AND_A28_B31, A[28], B[31]);
    wire P_A28_B31, Cout_A28_B31;
    full_adder add_a28_b31(P_A28_B31, Cout_A28_B31, P_A29_B30, AND_A28_B31, Cout_A28_B30);

    wire AND_A29_B31;
    nand and_a29_b31(AND_A29_B31, A[29], B[31]);
    wire P_A29_B31, Cout_A29_B31;
    full_adder add_a29_b31(P_A29_B31, Cout_A29_B31, P_A30_B30, AND_A29_B31, Cout_A29_B30);

    wire AND_A30_B31;
    nand and_a30_b31(AND_A30_B31, A[30], B[31]);
    wire P_A30_B31, Cout_A30_B31;
    full_adder add_a30_b31(P_A30_B31, Cout_A30_B31, P_A31_B30, AND_A30_B31, Cout_A30_B30);

    wire AND_A31_B31;
    and and_a31_b31(AND_A31_B31, A[31], B[31]);
    wire P_A31_B31, Cout_A31_B31;
    half_adder add_a31_b31(P_A31_B31, Cout_A31_B31, AND_A31_B31, Cout_A31_B30);






    wire S_A0_B31, Cout_A0_B31_final;
    half_adder s_a0_b31(S_A0_B31, Cout_A0_B31_final, P_A1_B31, Cout_A0_B31);
    
    wire S_A1_B31, Cout_A1_B31_final;
    full_adder s_a1_b31(S_A1_B31, Cout_A1_B31_final, P_A2_B31, Cout_A1_B31, Cout_A0_B31_final);

    wire S_A2_B31, Cout_A2_B31_final;
    full_adder s_a2_b31(S_A2_B31, Cout_A2_B31_final, P_A3_B31, Cout_A2_B31, Cout_A1_B31_final);
    wire S_A3_B31, Cout_A3_B31_final;
    full_adder s_a3_b31(S_A3_B31, Cout_A3_B31_final, P_A4_B31, Cout_A3_B31, Cout_A2_B31_final);
    wire S_A4_B31, Cout_A4_B31_final;
    full_adder s_a4_b31(S_A4_B31, Cout_A4_B31_final, P_A5_B31, Cout_A4_B31, Cout_A3_B31_final);
    wire S_A5_B31, Cout_A5_B31_final;
    full_adder s_a5_b31(S_A5_B31, Cout_A5_B31_final, P_A6_B31, Cout_A5_B31, Cout_A4_B31_final);
    wire S_A6_B31, Cout_A6_B31_final;
    full_adder s_a6_b31(S_A6_B31, Cout_A6_B31_final, P_A7_B31, Cout_A6_B31, Cout_A5_B31_final);
    wire S_A7_B31, Cout_A7_B31_final;
    full_adder s_a7_b31(S_A7_B31, Cout_A7_B31_final, P_A8_B31, Cout_A7_B31, Cout_A6_B31_final);
    wire S_A8_B31, Cout_A8_B31_final;
    full_adder s_a8_b31(S_A8_B31, Cout_A8_B31_final, P_A9_B31, Cout_A8_B31, Cout_A7_B31_final);
    wire S_A9_B31, Cout_A9_B31_final;
    full_adder s_a9_b31(S_A9_B31, Cout_A9_B31_final, P_A10_B31, Cout_A9_B31, Cout_A8_B31_final);
    wire S_A10_B31, Cout_A10_B31_final;
    full_adder s_a10_b31(S_A10_B31, Cout_A10_B31_final, P_A11_B31, Cout_A10_B31, Cout_A9_B31_final);
    wire S_A11_B31, Cout_A11_B31_final;
    full_adder s_a11_b31(S_A11_B31, Cout_A11_B31_final, P_A12_B31, Cout_A11_B31, Cout_A10_B31_final);
    wire S_A12_B31, Cout_A12_B31_final;
    full_adder s_a12_b31(S_A12_B31, Cout_A12_B31_final, P_A13_B31, Cout_A12_B31, Cout_A11_B31_final);
    wire S_A13_B31, Cout_A13_B31_final;
    full_adder s_a13_b31(S_A13_B31, Cout_A13_B31_final, P_A14_B31, Cout_A13_B31, Cout_A12_B31_final);
    wire S_A14_B31, Cout_A14_B31_final;
    full_adder s_a14_b31(S_A14_B31, Cout_A14_B31_final, P_A15_B31, Cout_A14_B31, Cout_A13_B31_final);
    wire S_A15_B31, Cout_A15_B31_final;
    full_adder s_a15_b31(S_A15_B31, Cout_A15_B31_final, P_A16_B31, Cout_A15_B31, Cout_A14_B31_final);
    wire S_A16_B31, Cout_A16_B31_final;
    full_adder s_a16_b31(S_A16_B31, Cout_A16_B31_final, P_A17_B31, Cout_A16_B31, Cout_A15_B31_final);
    wire S_A17_B31, Cout_A17_B31_final;
    full_adder s_a17_b31(S_A17_B31, Cout_A17_B31_final, P_A18_B31, Cout_A17_B31, Cout_A16_B31_final);
    wire S_A18_B31, Cout_A18_B31_final;
    full_adder s_a18_b31(S_A18_B31, Cout_A18_B31_final, P_A19_B31, Cout_A18_B31, Cout_A17_B31_final);
    wire S_A19_B31, Cout_A19_B31_final;
    full_adder s_a19_b31(S_A19_B31, Cout_A19_B31_final, P_A20_B31, Cout_A19_B31, Cout_A18_B31_final);
    wire S_A20_B31, Cout_A20_B31_final;
    full_adder s_a20_b31(S_A20_B31, Cout_A20_B31_final, P_A21_B31, Cout_A20_B31, Cout_A19_B31_final);
    wire S_A21_B31, Cout_A21_B31_final;
    full_adder s_a21_b31(S_A21_B31, Cout_A21_B31_final, P_A22_B31, Cout_A21_B31, Cout_A20_B31_final);
    wire S_A22_B31, Cout_A22_B31_final;
    full_adder s_a22_b31(S_A22_B31, Cout_A22_B31_final, P_A23_B31, Cout_A22_B31, Cout_A21_B31_final);
    wire S_A23_B31, Cout_A23_B31_final;
    full_adder s_a23_b31(S_A23_B31, Cout_A23_B31_final, P_A24_B31, Cout_A23_B31, Cout_A22_B31_final);
    wire S_A24_B31, Cout_A24_B31_final;
    full_adder s_a24_b31(S_A24_B31, Cout_A24_B31_final, P_A25_B31, Cout_A24_B31, Cout_A23_B31_final);
    wire S_A25_B31, Cout_A25_B31_final;
    full_adder s_a25_b31(S_A25_B31, Cout_A25_B31_final, P_A26_B31, Cout_A25_B31, Cout_A24_B31_final);
    wire S_A26_B31, Cout_A26_B31_final;
    full_adder s_a26_b31(S_A26_B31, Cout_A26_B31_final, P_A27_B31, Cout_A26_B31, Cout_A25_B31_final);
    wire S_A27_B31, Cout_A27_B31_final;
    full_adder s_a27_b31(S_A27_B31, Cout_A27_B31_final, P_A28_B31, Cout_A27_B31, Cout_A26_B31_final);
    wire S_A28_B31, Cout_A28_B31_final;
    full_adder s_a28_b31(S_A28_B31, Cout_A28_B31_final, P_A29_B31, Cout_A28_B31, Cout_A27_B31_final);
    wire S_A29_B31, Cout_A29_B31_final;
    full_adder s_a29_b31(S_A29_B31, Cout_A29_B31_final, P_A30_B31, Cout_A29_B31, Cout_A28_B31_final);
    wire S_A30_B31, Cout_A30_B31_final;
    full_adder s_a30_b31(S_A30_B31, Cout_A30_B31_final, P_A31_B31, Cout_A30_B31, Cout_A29_B31_final);
    wire S_A31_B31, Cout_A31_B31_final;
    full_adder s_a31_b31(S_A31_B31, Cout_A31_B31_final, single_one, Cout_A31_B31, Cout_A30_B31_final);

    


    assign P[0] = P_A0_B0;
    assign P[1] = P_A0_B1;
    assign P[2] = P_A0_B2;
    assign P[3] = P_A0_B3;
    assign P[4] = P_A0_B4;
    assign P[5] = P_A0_B5;
    assign P[6] = P_A0_B6;
    assign P[7] = P_A0_B7;
    assign P[8] = P_A0_B8;
    assign P[9] = P_A0_B9;
    assign P[10] =  P_A0_B10;
    assign P[11] =  P_A0_B11;
    assign P[12] =  P_A0_B12;
    assign P[13] =  P_A0_B13;
    assign P[14] =  P_A0_B14;
    assign P[15] =  P_A0_B15;
    assign P[16] =  P_A0_B16;
    assign P[17] =  P_A0_B17;
    assign P[18] =  P_A0_B18;
    assign P[19] =  P_A0_B19;
    assign P[20] =  P_A0_B20;
    assign P[21] =  P_A0_B21;
    assign P[22] =  P_A0_B22;
    assign P[23] =  P_A0_B23;
    assign P[24] =  P_A0_B24;
    assign P[25] =  P_A0_B25;
    assign P[26] =  P_A0_B26;
    assign P[27] =  P_A0_B27;
    assign P[28] =  P_A0_B28;
    assign P[29] =  P_A0_B29;
    assign P[30] =  P_A0_B30;
    assign P[31] =  P_A0_B31;

    assign P[32] = S_A0_B31;
    assign P[33] = S_A1_B31;
    assign P[34] = S_A2_B31;
    assign P[35] = S_A3_B31;
    assign P[36] = S_A4_B31;
    assign P[37] = S_A5_B31;
    assign P[38] = S_A6_B31;
    assign P[39] = S_A7_B31;
    assign P[40] = S_A8_B31;
    assign P[41] = S_A9_B31;
    assign P[42] = S_A10_B31;
    assign P[43] = S_A11_B31;
    assign P[44] = S_A12_B31;
    assign P[45] = S_A13_B31;
    assign P[46] = S_A14_B31;
    assign P[47] = S_A15_B31;
    assign P[48] = S_A16_B31;
    assign P[49] = S_A17_B31;
    assign P[50] = S_A18_B31;
    assign P[51] = S_A19_B31;
    assign P[52] = S_A20_B31;
    assign P[53] = S_A21_B31;
    assign P[54] = S_A22_B31;
    assign P[55] = S_A23_B31;
    assign P[56] = S_A24_B31;
    assign P[57] = S_A25_B31;
    assign P[58] = S_A26_B31;
    assign P[59] = S_A27_B31;
    assign P[60] = S_A28_B31;
    assign P[61] = S_A29_B31;
    assign P[62] = S_A30_B31;
    assign P[63] = S_A31_B31;    

    assign Pout[31:0] = P[31:0];

    wire [31:0] top32;
    assign top32[31:0] = P[63:32];

    assign ready = !zero;

    
    wire or_upper;
    assign or_upper = (P[63] | P[62] | P[61] | P[60] | P[59] | P[58] | P[57] | P[56] | P[55] | P[54] | P[53] | P[52] | P[51] | P[50] | P[49] | P[48] | P[47] | P[46] | P[45] | P[44] | P[43] | P[42] | P[41] | P[40] | P[39] | P[38] | P[37] | P[36] | P[35] | P[34] | P[33] | P[32]);
    
    wire and_upper;
    assign and_upper = (P[63] & P[62] & P[61] & P[60] & P[59] & P[58] & P[57] & P[56] & P[55] & P[54] & P[53] & P[52] & P[51] & P[50] & P[49] & P[48] & P[47] & P[46] & P[45] & P[44] & P[43] & P[42] & P[41] & P[40] & P[39] & P[38] & P[37] & P[36] & P[35] & P[34] & P[33] & P[32]);

    wire upper_ovf;
    assign upper_ovf = ~(and_upper | ~(or_upper));

    wire pos_a, pos_b, pos_p;
    assign pos_a = ~(A[31]);
    assign pos_b = ~(B[31]);
    assign pos_p = ~(P[31]);

    wire sign_ovf, s1, s2, s3, s4, s5;
    assign s1 = pos_a & pos_b & P[31];
    assign s2 = pos_a & B[31] & pos_p;
    assign s3 = A[31] & pos_b & pos_p;
    assign s4 = A[31] & B[31] & P[31];
    assign s5 = pos_a & pos_b & or_upper;
    assign sign_ovf = s1 | s2 | s3 | s4 | s5;

    assign Cout = upper_ovf | (sign_ovf & ~(a_zero | b_zero));


    // a or b is zero
    wire a_zero;
    assign a_zero = ~(A[31] | A[30] | A[29] | A[28] | A[27] | A[26] | A[25] | A[24] | A[23] | A[22] | A[21] | A[20] | A[19] | A[18] | A[17] | A[16] | A[15] | A[14] | A[13] | A[12] | A[11] | A[10] | A[9] | A[8] | A[7] | A[6] | A[5] | A[4] | A[3] | A[2] | A[1] | A[0]);
   
    wire b_zero;
    assign b_zero = ~(B[31] | B[30] | B[29] | B[28] | B[27] | B[26] | B[25] | B[24] | B[23] | B[22] | B[21] | B[20] | B[19] | B[18] | B[17] | B[16] | B[15] | B[14] | B[13] | B[12] | B[11] | B[10] | B[9] | B[8] | B[7] | B[6] | B[5] | B[4] | B[3] | B[2] | B[1] | B[0]);
   
    
    

endmodule